------------------------------------------------------------------------
-- Title      : Package for the clock_cross_pack logic
-- Project    : Tri-Mode Ethernet FIFO
------------------------------------------------------------------------
-- File       : clock_cross_pack.vhd
-- Author     : Xilinx Inc.
------------------------------------------------------------------------
-- (c) Copyright 2012 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
------------------------------------------------------------------------
-- Description:  This package contains all component declarations for
--               the entiries which make up the clock domain crossing
--               logic
------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

package clock_cross_pack is

  component sync_reset
  generic (
    DEPTH      : integer := 5
  );
  port (
    ARESET_IN  : in  std_logic;
    CLK        : in  std_logic;
    CE         : in  std_logic;
    SRESET_IN  : in  std_logic;
    RESET_OUT  : out std_logic
    );
  end component;

  component sync_block
  generic (
    INITIALISE : bit := '0';
    DEPTH      : integer := 5
  );
  port(
    clk        : in std_logic;
    reset      : in std_logic;
    data_in    : in std_logic;
    data_out   : out std_logic
  );
  end component;

  component bus_clk_cross
  generic (
    C_BUS_WIDTH    : integer range 2 to 64 := 8
  );
  port    (
    Clk_A_BUS_IN      : in  std_logic_vector(C_BUS_WIDTH-1 downto 0);    --  Clk A Bus In
    Clk_B             : in  std_logic;                                   --  Clk B
    Clk_B_Rst         : in  std_logic;                                   --  Clk B Reset
    stable_for_sample : in std_logic;
    ClkBBusOut     : out std_logic_vector(C_BUS_WIDTH-1 downto 0)     --  Clk B Bus Out
  );
  end component;

  component bus_and_enable_clk_cross
  generic (
    C_BUS_WIDTH    : integer range 2 to 64 := 8
  );
  port(
    ClkA          : in  std_logic;                                    --  Clk A Imput
    ClkA_EN       : in  std_logic;                                    --  Clk A Enable Input
    ClkARst       : in  std_logic;                                    --  Clk A Reset Input
    ClkASignalIn  : in  std_logic;                                    --  Clk A Signal In
    ClkABusIn     : in  std_logic_vector(C_BUS_WIDTH-1 downto 0);     --  Clk A Bus in
    ClkB          : in  std_logic;                                    --  Clk B Imput
    ClkB_EN       : in  std_logic;                                    --  Clk B Enable Input
    ClkBRst       : in  std_logic;                                    --  Clk B Reset Input
    ClkBSignalOut : out std_logic;                                    --  Clk B Signal Out
    ClkBBusOut    : out std_logic_vector(C_BUS_WIDTH-1 downto 0)      --  Clk B Bus Out
  );
  end component;

  component actv_hi_reset_clk_cross
  port    (
           ClkA               : in  std_logic;  --  Clock A input
           ClkAEN             : in  std_logic;  --  Enable signal clocked from clock A input
           ClkARst            : in  std_logic;  --  Clock A reset
           ClkAOutOfClkBRst   : out std_logic;  --  Held high until Clk B rst transitions LOW and is recognized by ClkA/CLKAEn
           ClkACombinedRstOut : out std_logic;  --  Held High until ClkBRst is detected LOW by ClkA/ClkAEn
           ClkB               : in  std_logic;  --  Clock B input
           ClkBEN             : in  std_logic;  --  Enable signal clocked from clock B input
           ClkBRst            : in  std_logic;  --  Clock B reset
           ClkBOutOfClkARst   : out std_logic;  --  Held high until Clk A rst transitions LOW and is recognized by ClkB/CLKBEn
           ClkBCombinedRstOut : out std_logic   --  Held High until ClkARst is detected LOW by ClkB/ClkBEn
          );
  end component;

  component actv_hi_pulse_clk_cross
  port    (
           ClkA          : in  std_logic; --  Clock A input
           ClkARst       : in  std_logic; --  Clock A reset
           ClkASignalIn  : in  std_logic; --  Signal clocked from Clock A input
           ClkB          : in  std_logic; --  Clock B input
           ClkBRst       : in  std_logic; --  Clock B reset
           ClkBSignalOut : out std_logic  --  Signal clocked from Clock B outout
          );
  end component;

end clock_cross_pack;


------------------------------------------------------------------------
-- Title      : CDC Sync Block (Synchroniser flip-flop pair)
-- Project    : AXI Ethernet Buffer
-------------------------------------------------------------------------------
-- File       : sync_block.vhd
-- Author     : Xilinx Inc.
--------------------------------------------------------------------------------
-- (c) Copyright 2001-2008 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Description: Used on signals crossing from one clock domain to another, this
--              is a multiple flip-flop pipeline, with all flops placed together
--              into the same slice.  Thus the routing delay between the two is
--              minimum to safe-guard against metastability issues.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library unisim;
use unisim.vcomponents.all;

entity sync_block is

  generic (
    INITIALISE : bit := '0';
    DEPTH      : integer := 5
  );

  port(
    clk        : in std_logic;
    reset      : in std_logic;
    data_in    : in std_logic;
    data_out   : out std_logic
  );

end sync_block;



architecture structural of sync_block is


  -- Internal Signals
  signal data_sync0 : std_logic;
  signal data_sync1 : std_logic;
  signal data_sync2 : std_logic;
  signal data_sync3 : std_logic;
  signal data_sync4 : std_logic;
  signal data_sync5 : std_logic;
  signal data_sync6 : std_logic;
  signal data_sync7 : std_logic;

  -- These ATTRIBUTES will stop timing errors being reported in back annotated SDF simulation.
  attribute async_reg               : string;
  attribute async_reg of data_sync0_i : label is "true";
  attribute async_reg of data_sync1_i : label is "true";
  attribute async_reg of data_sync2_i : label is "true";
  attribute async_reg of data_sync3_i : label is "true";
  attribute async_reg of data_sync4_i : label is "true";
  attribute async_reg of data_sync5_i : label is "true";
  attribute async_reg of data_sync6_i : label is "true";
  attribute async_reg of data_sync7_i : label is "true";
  attribute shreg_extract           : string;
  attribute shreg_extract of data_sync0_i : label is "no";
  attribute shreg_extract of data_sync1_i : label is "no";
  attribute shreg_extract of data_sync2_i : label is "no";
  attribute shreg_extract of data_sync3_i : label is "no";
  attribute shreg_extract of data_sync4_i : label is "no";
  attribute shreg_extract of data_sync5_i : label is "no";
  attribute shreg_extract of data_sync6_i : label is "no";
  attribute shreg_extract of data_sync7_i : label is "no";

begin


  data_sync0_i : FDRE
  generic map (
    INIT => INITIALISE
  )
  port map (
    C    => clk,
    CE   => '1',
    R    => reset,
    D    => data_in,
    Q    => data_sync0
  );

  data_sync1_i : FDRE
  generic map (
    INIT => INITIALISE
  )
  port map (
    C    => clk,
    CE   => '1',
    R    => reset,
    D    => data_sync0,
    Q    => data_sync1
  );

  data_sync2_i : FDRE
  generic map (
    INIT => INITIALISE
  )
  port map (
    C    => clk,
    CE   => '1',
    R    => reset,
    D    => data_sync1,
    Q    => data_sync2
  );

  data_sync3_i : FDRE
  generic map (
    INIT => INITIALISE
  )
  port map (
    C    => clk,
    CE   => '1',
    R    => reset,
    D    => data_sync2,
    Q    => data_sync3
  );

  data_sync4_i : FDRE
  generic map (
    INIT => INITIALISE
  )
  port map (
    C    => clk,
    CE   => '1',
    R    => reset,
    D    => data_sync3,
    Q    => data_sync4
  );

  data_sync5_i : FDRE
  generic map (
    INIT => INITIALISE
  )
  port map (
    C    => clk,
    CE   => '1',
    R    => reset,
    D    => data_sync4,
    Q    => data_sync5
  );

  data_sync6_i : FDRE
  generic map (
    INIT => INITIALISE
  )
  port map (
    C    => clk,
    CE   => '1',
    R    => reset,
    D    => data_sync5,
    Q    => data_sync6
  );

  data_sync7_i : FDRE
  generic map (
    INIT => INITIALISE
  )
  port map (
    C    => clk,
    CE   => '1',
    R    => reset,
    D    => data_sync6,
    Q    => data_sync7
  );

  data_out <= data_sync7;


end structural;


------------------------------------------------------------------------
-- Title      : Reset quasi-synchroniser
-- Project    : AXI Ethernet Buffer
------------------------------------------------------------------------
-- File       : sync_reset.vhd
-- Author     : Xilinx Inc.
------------------------------------------------------------------------
-- (c) Copyright 2001-2008 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
------------------------------------------------------------------------
-- Description: This reset synchronizer was derived from:
--              http://www.xilinx.com/support/techxclusives/global-techX19.htm
--              It is used to generate a reset signal which has a falling edge
--              synchronous with CLK; this allows predictable reset recovery
--              even using the asynchronous reset pins of register primitives.
-------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity sync_reset is

  generic (
    DEPTH      : integer := 5
  );
  port (
    ARESET_IN  : in  std_logic;         -- Active high asynchronous reset
    CLK        : in  std_logic;         -- clock to be sync'ed to
    CE         : in  std_logic;
    SRESET_IN  : in  std_logic;         -- Active high synchronous reset
    RESET_OUT  : out std_logic          -- "Synchronised" reset signal
    );

end sync_reset;

-------------------------------------------------------------------------------

architecture rtl of sync_reset is
    signal async_rst0 : std_logic := '1';
    signal async_rst1 : std_logic := '1';
    signal async_rst2 : std_logic := '1';
    signal async_rst3 : std_logic := '1';
    signal async_rst4 : std_logic := '1';
    signal sync_rst0  : std_logic := '1';
    signal sync_rst1  : std_logic := '1';

    attribute async_reg : string;
    attribute async_reg of async_rst0 : signal is "true";
    attribute async_reg of async_rst1 : signal is "true";
    attribute async_reg of async_rst2 : signal is "true";
    attribute async_reg of async_rst3 : signal is "true";
    attribute async_reg of async_rst4 : signal is "true";
    attribute async_reg of sync_rst0  : signal is "true";
    attribute async_reg of sync_rst1  : signal is "true";

    attribute shreg_extract               : string;
    attribute shreg_extract of async_rst0 : signal is "no";
    attribute shreg_extract of async_rst1 : signal is "no";
    attribute shreg_extract of async_rst2 : signal is "no";
    attribute shreg_extract of async_rst3 : signal is "no";
    attribute shreg_extract of async_rst4 : signal is "no";
    attribute shreg_extract of sync_rst0  : signal is "no";
    attribute shreg_extract of sync_rst1  : signal is "no";

begin  -- rtl

  -- Synchroniser process. In this case, 2 registers should pack into 1 slices.
  -- first two flops are asynchronously reset - 2 stage to ensure the reset is present for a full cycle
    P_RESET : process (CLK, ARESET_IN)
    begin
        if (ARESET_IN = '1') then
            async_rst0     <= '1';
        elsif CLK'event and CLK = '1' then
            async_rst0     <= '0';
        end if;
    end process P_RESET;

    RESET_SYNC_I : process (CLK, ARESET_IN)
    begin
        if (ARESET_IN = '1') then
            async_rst1   <= '1';
            async_rst2   <= '1';
            async_rst3   <= '1';
            async_rst4   <= '1';
        elsif CLK'event and CLK = '1' then
            async_rst1   <= async_rst0;
            async_rst2   <= async_rst1;
            async_rst3   <= async_rst2;
            async_rst4   <= async_rst3;
        end if;
    end process RESET_SYNC_I;

  -- second two flops are synchronously reset - this is used for all later flops
  -- and should ensure the reset is fully synchronous
    P_RESET_SYNC0 : process (CLK)
    begin
        if CLK'event and CLK = '1' then
            if (async_rst4 = '1' or SRESET_IN = '1') then
                sync_rst0     <= '1';
            elsif CE = '1' then
                sync_rst0     <= '0';
            end if;
        end if;
    end process P_RESET_SYNC0;

    P_RESET_SYNC1 : process (CLK)
    begin
        if CLK'event and CLK = '1' then
            if (async_rst4 = '1' or SRESET_IN = '1') then
                sync_rst1     <= '1';
            elsif CE = '1' then
                sync_rst1     <= sync_rst0;
            end if;
        end if;
    end process P_RESET_SYNC1;

    RESET_OUT <= sync_rst1;

end rtl;


------------------------------------------------------------------------------
-- actv_hi_reset_clk_cross - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2009, 2010 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--
------------------------------------------------------------------------------
-- Filename:        actv_hi_reset_clk_cross.vhd
-- Version:         v1.00a
-- Description:     This module converts an active high pulse from one clock to
--                   the other clock domain ensuring a pulse is detected
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              actv_hi_reset_clk_cross.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:      MSH
-- History:
-- MSH  10/28/2009
--        -- Initial design
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.clock_cross_pack.all;

entity actv_hi_reset_clk_cross is
    port    (
             ClkA               : in  std_logic;  --  Clock A input
             ClkAEN             : in  std_logic;  --  Enable signal clocked from clock A input
             ClkARst            : in  std_logic;  --  Clock A reset
             ClkAOutOfClkBRst   : out std_logic;  --  Held high until Clk B rst transitions LOW and is recognized by ClkA/CLKAEn
             ClkACombinedRstOut : out std_logic;  --  Held High until ClkBRst is detected LOW by ClkA/ClkAEn
             ClkB               : in  std_logic;  --  Clock B input
             ClkBEN             : in  std_logic;  --  Enable signal clocked from clock B input
             ClkBRst            : in  std_logic;  --  Clock B reset
             ClkBOutOfClkARst   : out std_logic;  --  Held high until Clk A rst transitions LOW and is recognized by ClkB/CLKBEn
             ClkBCombinedRstOut : out std_logic   --  Held High until ClkARst is detected LOW by ClkB/ClkBEn
            );
end actv_hi_reset_clk_cross;

architecture imp of actv_hi_reset_clk_cross is

  signal ClkBRstInternal    : std_logic;
  signal ClkARstInternal    : std_logic;

begin

  -- Notes: I don't know why clock enables are needed, but without visibility 
  -- I am keeping them to preserve original behaviour as close as possible

  ClkA_reset_inst: sync_reset
  port map (
    ARESET_IN  => ClkBRst,
    CLK        => ClkA,
	CE         => ClkAEN,
    SRESET_IN  => ClkARst,
    RESET_OUT  => ClkARstInternal
  );
  ClkAOutOfClkBRst   <= ClkARstInternal;
  ClkACombinedRstOut <= ClkARstInternal;


  ClkB_reset_inst: sync_reset
  port map (
    ARESET_IN  => ClkARst,
    CLK        => ClkB,
	CE         => ClkBEN,
    SRESET_IN  => ClkBRst,
    RESET_OUT  => ClkBRstInternal
  );
  ClkBOutOfClkARst   <= ClkBRstInternal;
  ClkBCombinedRstOut <= ClkBRstInternal;

	
end imp;


------------------------------------------------------------------------------
-- bus_clk_cross - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2009, 2010 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--
------------------------------------------------------------------------------
-- Filename:        bus_clk_cross.vhd
-- Version:         v1.00a
-- Description:     This module converts an active high pulse from one clock to
--                   the other clock domain ensuring a pulse is detected
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              bus_clk_cross.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:      MSH
-- History:
-- MSH  02/01/2010
--        -- Initial design
-- MBR  01/30/2013
--        -- rewritten with better metastability tolerance
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.clock_cross_pack.all;

entity bus_clk_cross is
  generic (
    C_BUS_WIDTH    : integer range 2 to 64 := 8
  );
  port    (
    Clk_A_BUS_IN      : in  std_logic_vector(C_BUS_WIDTH-1 downto 0);    --  Clk A Bus In
    Clk_B             : in  std_logic;                                   --  Clk B
    Clk_B_Rst         : in  std_logic;                                   --  Clk B Reset
    stable_for_sample : in  std_logic;                                   --  synchronous to clkB but indicates that Clk_A_BUS_IN is stable
    ClkBBusOut     : out std_logic_vector(C_BUS_WIDTH-1 downto 0)     --  Clk B Bus Out
  );
end bus_clk_cross;

architecture imp of bus_clk_cross is

  signal ClkBAxiEthBClkCrsBusOut    : std_logic_vector(C_BUS_WIDTH-1 downto 0)  ; 
  attribute async_reg               : string;
  attribute async_reg of ClkBAxiEthBClkCrsBusOut : signal is "true";

begin

  ClkBBusOut <= ClkBAxiEthBClkCrsBusOut;

  REG_DATA_PROCESS : process (Clk_B)
  begin
      if (Clk_B'event and Clk_B = '1') then
        if (Clk_B_Rst = '1') then
          ClkBAxiEthBClkCrsBusOut   <= Clk_A_BUS_IN;
        elsif stable_for_sample = '1' then
          ClkBAxiEthBClkCrsBusOut   <= Clk_A_BUS_IN;
        end if;
      end if;
  end process;

end imp;


------------------------------------------------------------------------------
-- bus_and_enable_clk_cross - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2009, 2010 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--
------------------------------------------------------------------------------
-- Filename:        bus_and_enable_clk_cross.vhd
-- Version:         v1.00a
-- Description:     This module converts an active high pulse from one clock to
--                   the other clock domain ensuring a pulse is detected
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              bus_and_enable_clk_cross.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:      MW
-- History:
-- MW  05/17/2010
--        -- Initial design
-- MBR  01/29/2013
--        -- rewritten with better metastability tolerance
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.clock_cross_pack.all;

library unisim;
use unisim.vcomponents.all;


entity bus_and_enable_clk_cross is
  generic (
    C_BUS_WIDTH    : integer range 2 to 64 := 8
  );
  port(
    ClkA          : in  std_logic;                                    --  Clk A Imput
    ClkA_EN       : in  std_logic;                                    --  Clk A Enable Input
    ClkARst       : in  std_logic;                                    --  Clk A Reset Input
    ClkASignalIn  : in  std_logic;                                    --  Clk A Signal In
    ClkABusIn     : in  std_logic_vector(C_BUS_WIDTH-1 downto 0);     --  Clk A Bus in
    ClkB          : in  std_logic;                                    --  Clk B Imput
    ClkB_EN       : in  std_logic;                                    --  Clk B Enable Input
    ClkBRst       : in  std_logic;                                    --  Clk B Reset Input
    ClkBSignalOut : out std_logic;                                    --  Clk B Signal Out
    ClkBBusOut    : out std_logic_vector(C_BUS_WIDTH-1 downto 0)      --  Clk B Bus Out
  );
end bus_and_enable_clk_cross;


architecture imp of bus_and_enable_clk_cross is


  signal ClkASignalInReg         : std_logic;
  signal ClkASignalToggle        : std_logic := '0';
  signal ClkASignalToggleSync    : std_logic;
  signal ClkASignalToggleSyncReg : std_logic;
  signal clk_a2b_bus    : std_logic_vector(C_BUS_WIDTH-1 downto 0) := (others => '0');

  signal ClkBAxiEthBaEClkCrsBusOut    : std_logic_vector(C_BUS_WIDTH-1 downto 0) ;  
  attribute async_reg               : string;
  attribute async_reg of ClkBAxiEthBaEClkCrsBusOut : signal is "true";

begin

  ClkBBusOut <= ClkBAxiEthBaEClkCrsBusOut;

  -- Register pulse A
  process(ClkA)
  begin
    if rising_edge(ClkA) then
      if ClkARst = '1' then
        ClkASignalInReg  <= '0';
      elsif ClkA_EN = '1' then
        ClkASignalInReg <= ClkASignalIn;
      end if;
    end if;
  end process;


  -- Detect rising edge of pulse A and create a toggle
  process(ClkA)
  begin
      if rising_edge(ClkA) then
          if ClkARst = '1' then
              ClkASignalToggle <= '0';
              clk_a2b_bus      <= (others => '0');
          else
              if ClkA_EN = '1' then
                  if ClkASignalIn = '1' and ClkASignalInReg = '0' then
                      ClkASignalToggle <= not ClkASignalToggle;
                      clk_a2b_bus      <= ClkABusIn;
                  end if;
              end if;
          end if;
      end if;
  end process;


  -- Include the metastability synchroniser
  data_sync : sync_block
  port map (
    clk        => ClkB,
	reset      => ClkBRst,
    data_in    => ClkASignalToggle,
    data_out   => ClkASignalToggleSync
  );


  -- Create the pulse on clock domain B
  process(ClkB)
  begin
    if rising_edge(ClkB) then
      if ClkBRst = '1' then
        ClkASignalToggleSyncReg <= '0';
        ClkBSignalOut           <= '0';
      elsif ClkB_EN = '1' then
        ClkASignalToggleSyncReg <= ClkASignalToggleSync;
        ClkBSignalOut           <= ClkASignalToggleSync xor ClkASignalToggleSyncReg;
      end if;
    end if;
  end process;


  -- Sample the data on clock domain B
  process(ClkB)
  begin
    if rising_edge(ClkB) then
      if ClkBRst = '1' then
        ClkBAxiEthBaEClkCrsBusOut <= (others => '0');
      elsif ClkB_EN = '1' then
        if (ClkASignalToggleSync xor ClkASignalToggleSyncReg) = '1' then
          ClkBAxiEthBaEClkCrsBusOut <= clk_a2b_bus;
        end if;
      end if;
    end if;
  end process;


end imp;


------------------------------------------------------------------------------
-- actv_hi_pulse_clk_cross - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2009, 2010 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--
------------------------------------------------------------------------------
-- Filename:        actv_hi_pulse_clk_cross.vhd
-- Version:         v1.00a
-- Description:     This module converts an active high pulse from one clock to
--                   the other clock domain ensuring a pulse is detected
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              actv_hi_pulse_clk_cross.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:      MSH
-- History:
-- MSH  10/28/2009
--        -- Initial design
-- MBR  01/29/2013
--        -- rewritten with better metastability tolerance
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.clock_cross_pack.all;

library unisim;
use unisim.vcomponents.all;


entity actv_hi_pulse_clk_cross is
    port    (
             ClkA          : in  std_logic; --  Clock A input
             ClkARst       : in  std_logic; --  Clock A reset
             ClkASignalIn  : in  std_logic; --  Signal clocked from Clock A input
             ClkB          : in  std_logic; --  Clock B input
             ClkBRst       : in  std_logic; --  Clock B reset
             ClkBSignalOut : out std_logic  --  Signal clocked from Clock B outout
            );
end actv_hi_pulse_clk_cross;


architecture imp of actv_hi_pulse_clk_cross is


  signal ClkASignalInReg         : std_logic;
  signal ClkASignalToggle        : std_logic := '0';
  signal ClkASignalToggleSync    : std_logic;
  signal ClkASignalToggleSyncReg : std_logic;


begin


  -- Register pulse A
  process(ClkA)
  begin
    if rising_edge(ClkA) then
      if ClkARst = '1' then
        ClkASignalInReg  <= '0';
      else
        ClkASignalInReg <= ClkASignalIn;
      end if;
    end if;
  end process;


  -- Detect rising edge of pulse A and create a toggle
  process(ClkA)
  begin
      if rising_edge(ClkA) then
          if ClkARst = '1' then
              ClkASignalToggle <= '0';
          else
              if ClkASignalIn = '1' and ClkASignalInReg = '0' then
                  ClkASignalToggle <= not ClkASignalToggle;
              else
                  ClkASignalToggle <= ClkASignalToggle;
              end if;
          end if;
      end if;
  end process;


  -- Include the metastability synchroniser
  data_sync : sync_block
  port map (
    clk        => ClkB,
	reset      => ClkBRst,
    data_in    => ClkASignalToggle,
    data_out   => ClkASignalToggleSync
  );


  -- Create the pulse on clock domain B
  process(ClkB)
  begin
    if rising_edge(ClkB) then
      if ClkBRst = '1' then
        ClkASignalToggleSyncReg <= '0';
        ClkBSignalOut           <= '0';
      else
        ClkASignalToggleSyncReg <= ClkASignalToggleSync;
        ClkBSignalOut           <= ClkASignalToggleSync xor ClkASignalToggleSyncReg;
      end if;
    end if;
  end process;


end imp;


-------------------------------------------------------------------------------
-- basic_sfifo_fg.vhd
-------------------------------------------------------------------------------
--
-- *************************************************************************
--
-- (c) Copyright 2010-2011 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-- *************************************************************************
--
-------------------------------------------------------------------------------
-- Filename:        basic_sfifo_fg.vhd
--
-- Description:     
-- This HDL file implements a basic synchronous (single clock) fifo using the
-- FIFO Generator tool. It is intended to offer a simple interface to the user
-- with the complexity of the FIFO Generator interface hidden from the user.               
--                  
-- Note that in normal op mode (not First Word Fall Through FWFT) the data count
-- output goes to zero when the FIFO goes full. This the way FIFO Generator works.
--                 
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              basic_sfifo_fg.vhd
--                 |
--                 |-- fifo_generator_v13_2
--
-------------------------------------------------------------------------------
-- Revision History:
--
--
-- Author:          DET
-- Revision:        $Revision: 1.0 $
-- Date:            $3/07/2011$
--
-- History:
--   DET   3/07/2011       Initial Version
-- 
-------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


--library fifo_generator_v13_2;
--use fifo_generator_v13_2.all;

Library xpm;
use xpm.vcomponents.all;

-------------------------------------------------------------------------------
entity basic_sfifo_fg is
  generic (
    
    C_DWIDTH                      : Integer :=  32 ;
      -- FIFO data Width (Read and write data ports are symetric)
    
    C_DEPTH                       : Integer := 512 ;
      -- FIFO Depth (set to power of 2)
 
    C_HAS_DATA_COUNT              : integer :=   1 ;
      -- 0 = Data Count output not needed
      -- 1 = Data Count output needed 
    
    C_DATA_COUNT_WIDTH            : integer :=  10 ;
    -- Data Count bit width (Max value is log2(C_DEPTH))
 
    C_IMPLEMENTATION_TYPE         : integer range 0 to 1 := 0;  
      --  0 = Common Clock BRAM / Distributed RAM (Synchronous FIFO)
      --  1 = Common Clock Shift Register (Synchronous FIFO)
    
    C_MEMORY_TYPE                 : integer := 1;
      --   0 = Any
      --   1 = BRAM
      --   2 = Distributed Memory  
      --   3 = Shift Registers
 
    C_PRELOAD_REGS                : integer := 1; 
      -- 0 = normal
      -- 1 = FWFT            
    
    C_PRELOAD_LATENCY             : integer := 0;              
      -- 0 = FWFT            
      -- 1 = normal
    
    C_USE_FWFT_DATA_COUNT         : integer := 0; 
      -- 0 = normal            
      -- 1 for FWFT
    C_SYNCHRONIZER_STAGE          : integer := 2;   -- valid values are 0 to 8;
 
    C_FAMILY                      : string  := "virtex6"
  
    );
  port (
    CLK                           : IN  std_logic := '0';
    DIN                           : IN  std_logic_vector(C_DWIDTH-1 DOWNTO 0) := (OTHERS => '0');
    RD_EN                         : IN  std_logic := '0';  
    SRST                          : IN  std_logic := '0';
    WR_EN                         : IN  std_logic := '0';
    DATA_COUNT                    : OUT std_logic_vector(C_DATA_COUNT_WIDTH-1 DOWNTO 0);
    DOUT                          : OUT std_logic_vector(C_DWIDTH-1 DOWNTO 0);
    EMPTY                         : OUT std_logic;
    FULL                          : OUT std_logic
    );
end entity basic_sfifo_fg;


architecture implementation of basic_sfifo_fg is
 -- Function delarations 

function log2(x : natural) return integer is
  variable i  : integer := 0;
  variable val: integer := 1;
begin
  if x = 0 then return 0;
  else
    for j in 0 to 29 loop -- for loop for XST 
      if val >= x then null;
      else
        i := i+1;
        val := val*2;
      end if;
    end loop;
  -- synthesis translate_off
    assert val >= x
      report "Function log2 received argument larger" &
             " than its capability of 2^30. "
      severity failure;
  -- synthesis translate_on
    return i;
  end if;
end function log2;

  FUNCTION if_then_else (
    condition : BOOLEAN;
    true_case : STRING;
    false_case : STRING)
  RETURN STRING IS
  BEGIN
    IF NOT condition THEN
      RETURN false_case;
    ELSE
      RETURN true_case;
    END IF;
  END if_then_else;

  FUNCTION PF_THRESH (
    DEPTH : INTEGER;
    RD_MODE: INTEGER)
  RETURN INTEGER IS
      VARIABLE FULL_THRESH : INTEGER;
  BEGIN
      FULL_THRESH := (DEPTH-3)-(RD_MODE*2);
      RETURN FULL_THRESH;
  END PF_THRESH;

  FUNCTION PE_THRESH (
    RD_MODE: INTEGER)
  RETURN INTEGER IS
      VARIABLE EMPTY_THRESH : INTEGER;
  BEGIN
      EMPTY_THRESH := 3+(RD_MODE*2);
      RETURN EMPTY_THRESH;
  END PE_THRESH;

  CONSTANT  P_FIFO_MEMORY_TYPE : STRING     := if_then_else( (C_MEMORY_TYPE = 0) , "auto" , if_then_else( (C_MEMORY_TYPE = 1) , "block" , if_then_else( (C_MEMORY_TYPE = 2) , "distributed" , if_then_else( (C_MEMORY_TYPE = 3) , "distributed" ,"auto"))));
  CONSTANT  P_USE_FWFT_DATA_COUNT : STRING     := if_then_else( (C_USE_FWFT_DATA_COUNT = 0) , "std" , "fwft");

  CONSTANT PROG_FULL_THRESH : INTEGER :=  PF_THRESH(C_DEPTH,C_USE_FWFT_DATA_COUNT);
  CONSTANT PROG_EMPTY_THRESH : INTEGER :=  PE_THRESH(C_USE_FWFT_DATA_COUNT);



  -- Constant Declarations  ----------------------------------------------
    Constant POINTER_WIDTH : integer := log2(C_DEPTH);
    
    -- Constant zeros for programmable threshold inputs
    signal PROG_RDTHRESH_ZEROS : std_logic_vector(POINTER_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
    signal PROG_WRTHRESH_ZEROS : std_logic_vector(POINTER_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
    
 -- Signals

  --Signals added to fix MTI and XSIM issues caused by fix for VCS issues not to use "LIBRARY_SCAN = TRUE"
    signal ALMOST_FULL         : std_logic;                       
    signal WR_ACK              : std_logic;                            
    signal OVERFLOW            : std_logic;                            
    signal VALID               : std_logic;                            
    signal UNDERFLOW           : std_logic;                            
    signal ALMOST_EMPTY        : std_logic;
    signal RD_DATA_COUNT       : std_logic_vector(C_DATA_COUNT_WIDTH-1 downto 0);
    signal WR_DATA_COUNT       : std_logic_vector(C_DATA_COUNT_WIDTH-1 downto 0);
    signal PROG_FULL           : std_logic;                 
    signal PROG_EMPTY          : std_logic;                 
    signal SBITERR             : std_logic;                 
    signal DBITERR             : std_logic;                  
    signal WR_RST_BUSY         : std_logic;                  
    signal RD_RST_BUSY         : std_logic;                  
    signal S_AXI_AWREADY       : std_logic;
    signal S_AXI_WREADY        : std_logic;
    signal S_AXI_BID           : std_logic_vector(3 DOWNTO 0);
    signal S_AXI_BRESP         : std_logic_vector(2-1 DOWNTO 0);
    signal S_AXI_BUSER         : std_logic_vector(0 downto 0);
    signal S_AXI_BVALID        : std_logic;

    -- AXI Full/Lite Master Write Channel (Read side)
    signal M_AXI_AWID          : std_logic_vector(3 DOWNTO 0);
    signal M_AXI_AWADDR        : std_logic_vector(31 DOWNTO 0);
    signal M_AXI_AWLEN         : std_logic_vector(8-1 DOWNTO 0);
    signal M_AXI_AWSIZE        : std_logic_vector(3-1 DOWNTO 0);
    signal M_AXI_AWBURST       : std_logic_vector(2-1 DOWNTO 0);
    signal M_AXI_AWLOCK        : std_logic_vector(2-1 DOWNTO 0);
    signal M_AXI_AWCACHE       : std_logic_vector(4-1 DOWNTO 0);
    signal M_AXI_AWPROT        : std_logic_vector(3-1 DOWNTO 0);
    signal M_AXI_AWQOS         : std_logic_vector(4-1 DOWNTO 0);
    signal M_AXI_AWREGION      : std_logic_vector(4-1 DOWNTO 0);
    signal M_AXI_AWUSER        : std_logic_vector(0 downto 0);
    signal M_AXI_AWVALID       : std_logic;
    signal M_AXI_WID           : std_logic_vector(3 DOWNTO 0);
    signal M_AXI_WDATA         : std_logic_vector(63 DOWNTO 0);
    signal M_AXI_WSTRB         : std_logic_vector(7 DOWNTO 0);
    signal M_AXI_WLAST         : std_logic;
    signal M_AXI_WUSER         : std_logic_vector(0 downto 0);
    signal M_AXI_WVALID        : std_logic;
    signal M_AXI_BREADY        : std_logic;

    -- AXI Full/Lite Slave Read Channel (Write side)
    signal S_AXI_ARREADY       : std_logic;
    signal S_AXI_RID           : std_logic_vector(3 DOWNTO 0);       
    signal S_AXI_RDATA         : std_logic_vector(63 DOWNTO 0); 
    signal S_AXI_RRESP         : std_logic_vector(2-1 DOWNTO 0);
    signal S_AXI_RLAST         : std_logic;
    signal S_AXI_RUSER         : std_logic_vector(0 downto 0);
    signal S_AXI_RVALID        : std_logic;

    -- AXI Full/Lite Master Read Channel (Read side)
    signal M_AXI_ARID          : std_logic_vector(3 DOWNTO 0);        
    signal M_AXI_ARADDR        : std_logic_vector(31 DOWNTO 0);  
    signal M_AXI_ARLEN         : std_logic_vector(8-1 DOWNTO 0);
    signal M_AXI_ARSIZE        : std_logic_vector(3-1 DOWNTO 0);
    signal M_AXI_ARBURST       : std_logic_vector(2-1 DOWNTO 0);
    signal M_AXI_ARLOCK        : std_logic_vector(2-1 DOWNTO 0);
    signal M_AXI_ARCACHE       : std_logic_vector(4-1 DOWNTO 0);
    signal M_AXI_ARPROT        : std_logic_vector(3-1 DOWNTO 0);
    signal M_AXI_ARQOS         : std_logic_vector(4-1 DOWNTO 0);
    signal M_AXI_ARREGION      : std_logic_vector(4-1 DOWNTO 0);
    signal M_AXI_ARUSER        : std_logic_vector(0 downto 0);
    signal M_AXI_ARVALID       : std_logic;
    signal M_AXI_RREADY        : std_logic;

    -- AXI Streaming Slave Signals (Write side)
    signal S_AXIS_TREADY       : std_logic;

    -- AXI Streaming Master Signals (Read side)
    signal M_AXIS_TVALID       : std_logic;
    signal M_AXIS_TDATA        : std_logic_vector(63 DOWNTO 0);
    signal M_AXIS_TSTRB        : std_logic_vector(3 DOWNTO 0);
    signal M_AXIS_TKEEP        : std_logic_vector(3 DOWNTO 0);
    signal M_AXIS_TLAST        : std_logic;
    signal M_AXIS_TID          : std_logic_vector(7 DOWNTO 0);
    signal M_AXIS_TDEST        : std_logic_vector(3 DOWNTO 0);
    signal M_AXIS_TUSER        : std_logic_vector(3 DOWNTO 0);

    -- AXI Full/Lite Write Address Channel Signals
    signal AXI_AW_DATA_COUNT    : std_logic_vector(4 DOWNTO 0);
    signal AXI_AW_WR_DATA_COUNT : std_logic_vector(4 DOWNTO 0);
    signal AXI_AW_RD_DATA_COUNT : std_logic_vector(4 DOWNTO 0);
    signal AXI_AW_SBITERR       : std_logic;
    signal AXI_AW_DBITERR       : std_logic;
    signal AXI_AW_OVERFLOW      : std_logic;
    signal AXI_AW_UNDERFLOW     : std_logic;
    signal AXI_AW_PROG_FULL     : STD_LOGIC;
    signal AXI_AW_PROG_EMPTY    : STD_LOGIC;


    -- AXI Full/Lite Write Data Channel Signals
    signal AXI_W_DATA_COUNT     : std_logic_vector(10 DOWNTO 0);
    signal AXI_W_WR_DATA_COUNT  : std_logic_vector(10 DOWNTO 0);
    signal AXI_W_RD_DATA_COUNT  : std_logic_vector(10 DOWNTO 0);
    signal AXI_W_SBITERR        : std_logic;
    signal AXI_W_DBITERR        : std_logic;
    signal AXI_W_OVERFLOW       : std_logic;
    signal AXI_W_UNDERFLOW      : std_logic;
    signal AXI_W_PROG_FULL      : STD_LOGIC;
    signal AXI_W_PROG_EMPTY     : STD_LOGIC;

    -- AXI Full/Lite Write Response Channel Signals
    signal AXI_B_DATA_COUNT     : std_logic_vector(4 DOWNTO 0);
    signal AXI_B_WR_DATA_COUNT  : std_logic_vector(4 DOWNTO 0);
    signal AXI_B_RD_DATA_COUNT  : std_logic_vector(4 DOWNTO 0);
    signal AXI_B_SBITERR        : std_logic;
    signal AXI_B_DBITERR        : std_logic;
    signal AXI_B_OVERFLOW       : std_logic;
    signal AXI_B_UNDERFLOW      : std_logic;
    signal AXI_B_PROG_FULL      : STD_LOGIC;
    signal AXI_B_PROG_EMPTY     : STD_LOGIC;

    -- AXI Full/Lite Read Address Channel Signals
    signal AXI_AR_DATA_COUNT    : std_logic_vector(4 DOWNTO 0);
    signal AXI_AR_WR_DATA_COUNT : std_logic_vector(4 DOWNTO 0);
    signal AXI_AR_RD_DATA_COUNT : std_logic_vector(4 DOWNTO 0);
    signal AXI_AR_SBITERR       : std_logic;
    signal AXI_AR_DBITERR       : std_logic;
    signal AXI_AR_OVERFLOW      : std_logic;
    signal AXI_AR_UNDERFLOW     : std_logic;
    signal AXI_AR_PROG_FULL     : STD_LOGIC;
    signal AXI_AR_PROG_EMPTY    : STD_LOGIC;

    -- AXI Full/Lite Read Data Channel Signals
    signal AXI_R_DATA_COUNT     : std_logic_vector(10 DOWNTO 0);
    signal AXI_R_WR_DATA_COUNT  : std_logic_vector(10 DOWNTO 0);
    signal AXI_R_RD_DATA_COUNT  : std_logic_vector(10 DOWNTO 0);
    signal AXI_R_SBITERR        : std_logic;
    signal AXI_R_DBITERR        : std_logic;
    signal AXI_R_OVERFLOW       : std_logic;
    signal AXI_R_UNDERFLOW      : std_logic;
    signal AXI_R_PROG_FULL      : STD_LOGIC;
    signal AXI_R_PROG_EMPTY     : STD_LOGIC;

    -- AXI Streaming FIFO Related Signals
    signal AXIS_DATA_COUNT      : std_logic_vector(10 DOWNTO 0);
    signal AXIS_WR_DATA_COUNT   : std_logic_vector(10 DOWNTO 0);
    signal AXIS_RD_DATA_COUNT   : std_logic_vector(10 DOWNTO 0);
    signal AXIS_SBITERR         : std_logic;
    signal AXIS_DBITERR         : std_logic;
    signal AXIS_OVERFLOW        : std_logic;
    signal AXIS_UNDERFLOW       : std_logic;
    signal AXIS_PROG_FULL       : STD_LOGIC;
    signal AXIS_PROG_EMPTY      : STD_LOGIC;


begin --(architecture implementation)

 

  -------------------------------------------------------------------------------
  -- Instantiate the generalized FIFO Generator instance
  --
  -- NOTE:
  -- DO NOT CHANGE TO DIRECT ENTITY INSTANTIATION!!!
  -- This is a Coregen FIFO Generator Call module for 
  -- BRAM implementations of a basic Sync FIFO
  --
  -------------------------------------------------------------------------------
I_BASIC_SFIFO: xpm_fifo_sync
  generic map (

    FIFO_MEMORY_TYPE         => P_FIFO_MEMORY_TYPE,           --string; "auto", "block", "distributed", or "ultra" ;
    ECC_MODE                 => "no_ecc",         --string; "no_ecc" or "en_ecc";
    FIFO_WRITE_DEPTH         => C_DEPTH,             --positive integer
    WRITE_DATA_WIDTH         => C_DWIDTH,               --positive integer
    WR_DATA_COUNT_WIDTH      => C_DATA_COUNT_WIDTH,               --positive integer
    PROG_FULL_THRESH         => PROG_FULL_THRESH,               --positive integer
    FULL_RESET_VALUE         => 0,                --positive integer; 0 or 1;
    USE_ADV_FEATURES         => "0707",           --string; "0000" to "1F1F";
    READ_MODE                => P_USE_FWFT_DATA_COUNT,            --string; "std" or "fwft";
    FIFO_READ_LATENCY        => 1,                --positive integer;
    READ_DATA_WIDTH          => C_DWIDTH,               --positive integer
    RD_DATA_COUNT_WIDTH      => C_DATA_COUNT_WIDTH,               --positive integer
    PROG_EMPTY_THRESH        => PROG_EMPTY_THRESH,               --positive integer
    DOUT_RESET_VALUE         => "0",              --string
    WAKEUP_TIME              => 0                 --positive integer; 0 or 2;
  )
  port map (

    rst              => SRST,
    wr_clk           => CLK,
    wr_en            => WR_EN,
    din              => DIN,
    full             => FULL,
    overflow         => OVERFLOW,
    wr_rst_busy      => WR_RST_BUSY,
    prog_full        => PROG_FULL,
    wr_data_count    => DATA_COUNT,
    almost_full      => ALMOST_FULL,
    wr_ack           => WR_ACK,
    rd_en            => RD_EN,
    dout             => DOUT,
    empty            => EMPTY,
    underflow        => UNDERFLOW,
    rd_rst_busy      => RD_RST_BUSY,
    prog_empty       => PROG_EMPTY,
    rd_data_count    => RD_DATA_COUNT,
    almost_empty     => ALMOST_EMPTY,
    data_valid       => VALID,
    sleep            => '0',
    injectsbiterr    => '0',
    injectdbiterr    => '0',
    sbiterr          => SBITERR,
    dbiterr          => DBITERR
  );



--  I_BASIC_SFIFO : entity fifo_generator_v13_2.fifo_generator_v13_2 
--    generic map(
--      C_COMMON_CLOCK                 =>  1,                                           
--      C_COUNT_TYPE                   =>  0,                                           
--      C_DATA_COUNT_WIDTH             =>  C_DATA_COUNT_WIDTH,   
--      C_DEFAULT_VALUE                =>  "BlankString",        
--      C_DIN_WIDTH                    =>  C_DWIDTH,                          
--      C_DOUT_RST_VAL                 =>  "0",
--      C_DOUT_WIDTH                   =>  C_DWIDTH,
--      C_ENABLE_RLOCS                 =>  0,  -- n0
--      C_FAMILY                       =>  C_FAMILY,
--      C_HAS_ALMOST_EMPTY             =>  0,  -- n0
--      C_HAS_ALMOST_FULL              =>  0,  -- n0        
--      C_HAS_BACKUP                   =>  0,  -- n0 
--      C_HAS_DATA_COUNT               =>  C_HAS_DATA_COUNT,
--      C_HAS_MEMINIT_FILE             =>  0,  -- n0
--      C_HAS_OVERFLOW                 =>  0,  -- n0
--      C_HAS_RD_DATA_COUNT            =>  0,  -- n0
--      C_HAS_RD_RST                   =>  0,  -- n0
--      C_HAS_RST                      =>  0,  -- n0
--      C_HAS_SRST                     =>  1,  -- yes
--      C_HAS_UNDERFLOW                =>  0,  -- n0
--      C_HAS_VALID                    =>  0,  -- n0
--      C_HAS_WR_ACK                   =>  0,  -- n0
--      C_HAS_WR_DATA_COUNT            =>  0,  -- n0
--      C_HAS_WR_RST                   =>  0,  -- n0
--      C_IMPLEMENTATION_TYPE          =>  0,  -- Common clock BRAM
--      C_INIT_WR_PNTR_VAL             =>  0,
--      C_MEMORY_TYPE                  =>  C_MEMORY_TYPE,
--      C_MIF_FILE_NAME                =>  "BlankString",
--      C_OPTIMIZATION_MODE            =>  0,
--      C_OVERFLOW_LOW                 =>  0,
--      C_PRELOAD_LATENCY              =>  C_PRELOAD_LATENCY,                                        
--      C_PRELOAD_REGS                 =>  C_PRELOAD_REGS,                                    
--      C_PRIM_FIFO_TYPE               =>  "512x36",
--      C_PROG_EMPTY_THRESH_ASSERT_VAL =>  0,
--      C_PROG_EMPTY_THRESH_NEGATE_VAL =>  0,
--      C_PROG_EMPTY_TYPE              =>  0,
--      C_PROG_FULL_THRESH_ASSERT_VAL  =>  0,
--      C_PROG_FULL_THRESH_NEGATE_VAL  =>  0,
--      C_PROG_FULL_TYPE               =>  0,
--      C_RD_DATA_COUNT_WIDTH          =>  C_DATA_COUNT_WIDTH,
--      C_RD_DEPTH                     =>  C_DEPTH,
--      C_RD_FREQ                      =>  1,
--      C_RD_PNTR_WIDTH                =>  POINTER_WIDTH,
--      C_UNDERFLOW_LOW                =>  0,
--      C_USE_DOUT_RST                 =>  1,
--      C_USE_EMBEDDED_REG             =>  0,
--      C_USE_FIFO16_FLAGS             =>  0,
--      C_USE_FWFT_DATA_COUNT          =>  C_USE_FWFT_DATA_COUNT,
--      C_VALID_LOW                    =>  0,
--      C_WR_ACK_LOW                   =>  0,
--      C_WR_DATA_COUNT_WIDTH          =>  C_DATA_COUNT_WIDTH,
--      C_WR_DEPTH                     =>  C_DEPTH,
--      C_WR_FREQ                      =>  1,
--      C_WR_PNTR_WIDTH                =>  POINTER_WIDTH,
--      C_WR_RESPONSE_LATENCY          =>  1,
--      C_USE_ECC                      =>  0,
--      C_FULL_FLAGS_RST_VAL           =>  1,
--      C_ENABLE_RST_SYNC              =>  1,
--      C_ERROR_INJECTION_TYPE         =>  0,
--      C_SYNCHRONIZER_STAGE           =>  C_SYNCHRONIZER_STAGE,
--      C_HAS_INT_CLK                  =>  0,
--      C_MSGON_VAL                    =>  1,
--      
--
--      -- AXI Interface related parameters start here
--      C_INTERFACE_TYPE               =>  0,    --           : integer := 0; -- 0: Native Interface; 1: AXI Interface
--      C_AXI_TYPE                     =>  0,    --           : integer := 0; -- 0: AXI Stream; 1: AXI Full; 2: AXI Lite
--      C_HAS_AXI_WR_CHANNEL           =>  0,    --           : integer := 0;
--      C_HAS_AXI_RD_CHANNEL           =>  0,    --           : integer := 0;
--      C_HAS_SLAVE_CE                 =>  0,    --           : integer := 0;
--      C_HAS_MASTER_CE                =>  0,    --           : integer := 0;
--      C_ADD_NGC_CONSTRAINT           =>  0,    --           : integer := 0;
--      C_USE_COMMON_OVERFLOW          =>  0,    --           : integer := 0;
--      C_USE_COMMON_UNDERFLOW         =>  0,    --           : integer := 0;
--      C_USE_DEFAULT_SETTINGS         =>  0,    --           : integer := 0;
--
--      -- AXI Full/Lite
--      C_AXI_ID_WIDTH                 =>  4 ,    --           : integer := 0;
--      C_AXI_ADDR_WIDTH               =>  32,    --           : integer := 0;
--      C_AXI_DATA_WIDTH               =>  64,    --           : integer := 0;
--      C_AXI_LEN_WIDTH                =>  8,     --           : integer := 8;
--      C_AXI_LOCK_WIDTH               =>  2,     --           : integer := 2;
--      C_HAS_AXI_ID                   =>  0,     --           : integer := 0;
--      C_HAS_AXI_AWUSER               =>  0 ,    --           : integer := 0;
--      C_HAS_AXI_WUSER                =>  0 ,    --           : integer := 0;
--      C_HAS_AXI_BUSER                =>  0 ,    --           : integer := 0;
--      C_HAS_AXI_ARUSER               =>  0 ,    --           : integer := 0;
--      C_HAS_AXI_RUSER                =>  0 ,    --           : integer := 0;
--      C_AXI_ARUSER_WIDTH             =>  1 ,    --           : integer := 0;
--      C_AXI_AWUSER_WIDTH             =>  1 ,    --           : integer := 0;
--      C_AXI_WUSER_WIDTH              =>  1 ,    --           : integer := 0;
--      C_AXI_BUSER_WIDTH              =>  1 ,    --           : integer := 0;
--      C_AXI_RUSER_WIDTH              =>  1 ,    --           : integer := 0;
--                                         
--      -- AXI Streaming
--      C_HAS_AXIS_TDATA               =>  0 ,    --           : integer := 0;
--      C_HAS_AXIS_TID                 =>  0 ,    --           : integer := 0;
--      C_HAS_AXIS_TDEST               =>  0 ,    --           : integer := 0;
--      C_HAS_AXIS_TUSER               =>  0 ,    --           : integer := 0;
--      C_HAS_AXIS_TREADY              =>  1 ,    --           : integer := 0;
--      C_HAS_AXIS_TLAST               =>  0 ,    --           : integer := 0;
--      C_HAS_AXIS_TSTRB               =>  0 ,    --           : integer := 0;
--      C_HAS_AXIS_TKEEP               =>  0 ,    --           : integer := 0;
--      C_AXIS_TDATA_WIDTH             =>  64,    --           : integer := 1;
--      C_AXIS_TID_WIDTH               =>  8 ,    --           : integer := 1;
--      C_AXIS_TDEST_WIDTH             =>  4 ,    --           : integer := 1;
--      C_AXIS_TUSER_WIDTH             =>  4 ,    --           : integer := 1;
--      C_AXIS_TSTRB_WIDTH             =>  4 ,    --           : integer := 1;
--      C_AXIS_TKEEP_WIDTH             =>  4 ,    --           : integer := 1;
--
--      -- AXI Channel Type
--      -- WACH --> Write Address Channel
--      -- WDCH --> Write Data Channel
--      -- WRCH --> Write Response Channel
--      -- RACH --> Read Address Channel
--      -- RDCH --> Read Data Channel
--      -- AXIS --> AXI Streaming
--      C_WACH_TYPE                   =>  0,    --            : integer := 0; -- 0 = FIFO; 1 = Register Slice; 2 = Pass Through Logic
--      C_WDCH_TYPE                   =>  0,    --            : integer := 0; -- 0 = FIFO; 1 = Register Slice; 2 = Pass Through Logie
--      C_WRCH_TYPE                   =>  0,    --            : integer := 0; -- 0 = FIFO; 1 = Register Slice; 2 = Pass Through Logie
--      C_RACH_TYPE                   =>  0,    --            : integer := 0; -- 0 = FIFO; 1 = Register Slice; 2 = Pass Through Logie
--      C_RDCH_TYPE                   =>  0,    --            : integer := 0; -- 0 = FIFO; 1 = Register Slice; 2 = Pass Through Logie
--      C_AXIS_TYPE                   =>  0,    --            : integer := 0; -- 0 = FIFO; 1 = Register Slice; 2 = Pass Through Logie
--
--      -- AXI Implementation Type
--      -- 1 = Common Clock Block RAM FIFO
--      -- 2 = Common Clock Distributed RAM FIFO
--      -- 11 = Independent Clock Block RAM FIFO
--      -- 12 = Independent Clock Distributed RAM FIFO
--      C_IMPLEMENTATION_TYPE_WACH    =>  1,    --            : integer := 0;
--      C_IMPLEMENTATION_TYPE_WDCH    =>  1,    --            : integer := 0;
--      C_IMPLEMENTATION_TYPE_WRCH    =>  1,    --            : integer := 0;
--      C_IMPLEMENTATION_TYPE_RACH    =>  1,    --            : integer := 0;
--      C_IMPLEMENTATION_TYPE_RDCH    =>  1,    --            : integer := 0;
--      C_IMPLEMENTATION_TYPE_AXIS    =>  1,    --            : integer := 0;
--
--      -- AXI FIFO Type
--      -- 0 = Data FIFO
--      -- 1 = Packet FIFO
--      -- 2 = Low Latency Data FIFO
--      C_APPLICATION_TYPE_WACH      =>  0,    --             : integer := 0;
--      C_APPLICATION_TYPE_WDCH      =>  0,    --             : integer := 0;
--      C_APPLICATION_TYPE_WRCH      =>  0,    --             : integer := 0;
--      C_APPLICATION_TYPE_RACH      =>  0,    --             : integer := 0;
--      C_APPLICATION_TYPE_RDCH      =>  0,    --             : integer := 0;
--      C_APPLICATION_TYPE_AXIS      =>  0,    --             : integer := 0;
--
--      -- Enable ECC
--      -- 0 = ECC disabled
--      -- 1 = ECC enabled
--      C_USE_ECC_WACH               =>  0,    --             : integer := 0;
--      C_USE_ECC_WDCH               =>  0,    --             : integer := 0;
--      C_USE_ECC_WRCH               =>  0,    --             : integer := 0;
--      C_USE_ECC_RACH               =>  0,    --             : integer := 0;
--      C_USE_ECC_RDCH               =>  0,    --             : integer := 0;
--      C_USE_ECC_AXIS               =>  0,    --             : integer := 0;
--
--      -- ECC Error Injection Type
--      -- 0 = No Error Injection
--      -- 1 = Single Bit Error Injection
--      -- 2 = Double Bit Error Injection
--      -- 3 = Single Bit and Double Bit Error Injection
--      C_ERROR_INJECTION_TYPE_WACH  =>  0,    --             : integer := 0;
--      C_ERROR_INJECTION_TYPE_WDCH  =>  0,    --             : integer := 0;
--      C_ERROR_INJECTION_TYPE_WRCH  =>  0,    --             : integer := 0;
--      C_ERROR_INJECTION_TYPE_RACH  =>  0,    --             : integer := 0;
--      C_ERROR_INJECTION_TYPE_RDCH  =>  0,    --             : integer := 0;
--      C_ERROR_INJECTION_TYPE_AXIS  =>  0,    --             : integer := 0;
--
--      -- Input Data Width
--      -- Accumulation of all AXI input signal's width
--      C_DIN_WIDTH_WACH                    =>  32,    --      : integer := 1;
--      C_DIN_WIDTH_WDCH                    =>  64,    --      : integer := 1;
--      C_DIN_WIDTH_WRCH                    =>  2 ,    --      : integer := 1;
--      C_DIN_WIDTH_RACH                    =>  32,    --      : integer := 1;
--      C_DIN_WIDTH_RDCH                    =>  64,    --      : integer := 1;
--      C_DIN_WIDTH_AXIS                    =>  1 ,    --      : integer := 1;
--
--      C_WR_DEPTH_WACH                     =>  16  ,   --      : integer := 16;
--      C_WR_DEPTH_WDCH                     =>  1024,   --      : integer := 16;
--      C_WR_DEPTH_WRCH                     =>  16  ,   --      : integer := 16;
--      C_WR_DEPTH_RACH                     =>  16  ,   --      : integer := 16;
--      C_WR_DEPTH_RDCH                     =>  1024,   --      : integer := 16;
--      C_WR_DEPTH_AXIS                     =>  1024,   --      : integer := 16;
--
--      C_WR_PNTR_WIDTH_WACH                =>  4 ,    --      : integer := 4;
--      C_WR_PNTR_WIDTH_WDCH                =>  10,    --      : integer := 4;
--      C_WR_PNTR_WIDTH_WRCH                =>  4 ,    --      : integer := 4;
--      C_WR_PNTR_WIDTH_RACH                =>  4 ,    --      : integer := 4;
--      C_WR_PNTR_WIDTH_RDCH                =>  10,    --      : integer := 4;
--      C_WR_PNTR_WIDTH_AXIS                =>  10,    --      : integer := 4;
--
--      C_HAS_DATA_COUNTS_WACH              =>  0,    --      : integer := 0;
--      C_HAS_DATA_COUNTS_WDCH              =>  0,    --      : integer := 0;
--      C_HAS_DATA_COUNTS_WRCH              =>  0,    --      : integer := 0;
--      C_HAS_DATA_COUNTS_RACH              =>  0,    --      : integer := 0;
--      C_HAS_DATA_COUNTS_RDCH              =>  0,    --      : integer := 0;
--      C_HAS_DATA_COUNTS_AXIS              =>  0,    --      : integer := 0;
--
--      C_HAS_PROG_FLAGS_WACH               =>  0,    --      : integer := 0;
--      C_HAS_PROG_FLAGS_WDCH               =>  0,    --      : integer := 0;
--      C_HAS_PROG_FLAGS_WRCH               =>  0,    --      : integer := 0;
--      C_HAS_PROG_FLAGS_RACH               =>  0,    --      : integer := 0;
--      C_HAS_PROG_FLAGS_RDCH               =>  0,    --      : integer := 0;
--      C_HAS_PROG_FLAGS_AXIS               =>  0,    --      : integer := 0;
--
--      C_PROG_FULL_TYPE_WACH               =>  5   ,    --      : integer := 0;
--      C_PROG_FULL_TYPE_WDCH               =>  5   ,    --      : integer := 0;
--      C_PROG_FULL_TYPE_WRCH               =>  5   ,    --      : integer := 0;
--      C_PROG_FULL_TYPE_RACH               =>  5   ,    --      : integer := 0;
--      C_PROG_FULL_TYPE_RDCH               =>  5   ,    --      : integer := 0;
--      C_PROG_FULL_TYPE_AXIS               =>  5   ,    --      : integer := 0;
--      C_PROG_FULL_THRESH_ASSERT_VAL_WACH  =>  1023,    --      : integer := 0;
--      C_PROG_FULL_THRESH_ASSERT_VAL_WDCH  =>  1023,    --      : integer := 0;
--      C_PROG_FULL_THRESH_ASSERT_VAL_WRCH  =>  1023,    --      : integer := 0;
--      C_PROG_FULL_THRESH_ASSERT_VAL_RACH  =>  1023,    --      : integer := 0;
--      C_PROG_FULL_THRESH_ASSERT_VAL_RDCH  =>  1023,    --      : integer := 0;
--      C_PROG_FULL_THRESH_ASSERT_VAL_AXIS  =>  1023,    --      : integer := 0;
--
--      C_PROG_EMPTY_TYPE_WACH              =>  5   ,    --      : integer := 0;
--      C_PROG_EMPTY_TYPE_WDCH              =>  5   ,    --      : integer := 0;
--      C_PROG_EMPTY_TYPE_WRCH              =>  5   ,    --      : integer := 0;
--      C_PROG_EMPTY_TYPE_RACH              =>  5   ,    --      : integer := 0;
--      C_PROG_EMPTY_TYPE_RDCH              =>  5   ,    --      : integer := 0;
--      C_PROG_EMPTY_TYPE_AXIS              =>  5   ,    --      : integer := 0;
--      C_PROG_EMPTY_THRESH_ASSERT_VAL_WACH =>  1022,    --      : integer := 0;
--      C_PROG_EMPTY_THRESH_ASSERT_VAL_WDCH =>  1022,    --      : integer := 0;
--      C_PROG_EMPTY_THRESH_ASSERT_VAL_WRCH =>  1022,    --      : integer := 0;
--      C_PROG_EMPTY_THRESH_ASSERT_VAL_RACH =>  1022,    --      : integer := 0;
--      C_PROG_EMPTY_THRESH_ASSERT_VAL_RDCH =>  1022,    --      : integer := 0;
--      C_PROG_EMPTY_THRESH_ASSERT_VAL_AXIS =>  1022,    --      : integer := 0;
--
--      C_REG_SLICE_MODE_WACH               =>  0,    --      : integer := 0;
--      C_REG_SLICE_MODE_WDCH               =>  0,    --      : integer := 0;
--      C_REG_SLICE_MODE_WRCH               =>  0,    --      : integer := 0;
--      C_REG_SLICE_MODE_RACH               =>  0,    --      : integer := 0;
--      C_REG_SLICE_MODE_RDCH               =>  0,    --      : integer := 0;
--      C_REG_SLICE_MODE_AXIS               =>  0     --      : integer := 0
--
--      )
--    port map(
--      backup                    =>  '0',                  
--      backup_marker             =>  '0',                  
--      clk                       =>  CLK,                  
--      rst                       =>  '0',                  
--      srst                      =>  SRST,          
--      wr_clk                    =>  '0',                  
--      wr_rst                    =>  '0',                  
--      rd_clk                    =>  '0',                  
--      rd_rst                    =>  '0',                  
--      din                       =>  DIN,                 -- uses this one            
--      wr_en                     =>  WR_EN,               -- uses this one            
--      rd_en                     =>  RD_EN,               -- uses this one            
--      prog_empty_thresh         =>  PROG_RDTHRESH_ZEROS,  
--      prog_empty_thresh_assert  =>  PROG_RDTHRESH_ZEROS,  
--      prog_empty_thresh_negate  =>  PROG_RDTHRESH_ZEROS,  
--      prog_full_thresh          =>  PROG_WRTHRESH_ZEROS,  
--      prog_full_thresh_assert   =>  PROG_WRTHRESH_ZEROS,  
--      prog_full_thresh_negate   =>  PROG_WRTHRESH_ZEROS,  
--      int_clk                   =>  '0',                  
--      injectdbiterr             =>  '0', 
--      injectsbiterr             =>  '0', 
--      sleep                     =>  '0',
--                                                                                                                             
--      dout                      =>  DOUT,                -- uses this one           
--      full                      =>  FULL,                -- uses this one           
--      almost_full               =>  ALMOST_FULL,                       
--      wr_ack                    =>  WR_ACK,                            
--      overflow                  =>  OVERFLOW,                            
--      empty                     =>  EMPTY,               -- uses this one
--      almost_empty              =>  ALMOST_EMPTY,                              
--      valid                     =>  VALID,                            
--      underflow                 =>  UNDERFLOW,                            
--      data_count                =>  DATA_COUNT,          -- uses this one          
--      rd_data_count             =>  RD_DATA_COUNT,                              
--      wr_data_count             =>  WR_DATA_COUNT,                              
--      prog_full                 =>  PROG_FULL,                              
--      prog_empty                =>  PROG_EMPTY,                              
--      sbiterr                   =>  SBITERR,                              
--      dbiterr                   =>  DBITERR,
--      wr_rst_busy               =>  WR_RST_BUSY,
--      rd_rst_busy               =>  RD_RST_BUSY,           
--
--      -- AXI Global Signal
--      m_aclk                    =>  '0',                   --       : IN  std_logic := '0';
--      s_aclk                    =>  '0',                   --       : IN  std_logic := '0';
--      s_aresetn                 =>  '0',                   --       : IN  std_logic := '0';
--      m_aclk_en                 =>  '0',                   --       : IN  std_logic := '0';
--      s_aclk_en                 =>  '0',                   --       : IN  std_logic := '0';
--
--      -- AXI Full/Lite Slave Write Channel (write side)
--      s_axi_awid                =>  "0000",         --(others => '0'),      --      : IN  std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awaddr              =>  "00000000000000000000000000000000",   --(others => '0'),      --      : IN  std_logic_vector(C_AXI_ADDR_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awlen               =>  "00000000",          --(others => '0'),      --      : IN  std_logic_vector(8-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awsize              =>  "000",          --(others => '0'),      --      : IN  std_logic_vector(3-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awburst             =>  "00",           --(others => '0'),      --      : IN  std_logic_vector(2-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awlock              =>  "00",           --(others => '0'),      --      : IN  std_logic_vector(2-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awcache             =>  "0000",         --(others => '0'),      --      : IN  std_logic_vector(4-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awprot              =>  "000",          --(others => '0'),      --      : IN  std_logic_vector(3-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awqos               =>  "0000",         --(others => '0'),      --      : IN  std_logic_vector(4-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awregion            =>  "0000",         --(others => '0'),      --      : IN  std_logic_vector(4-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awuser              =>  "0",            --(others => '0'),      --      : IN  std_logic_vector(C_AXI_AWUSER_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_awvalid             =>  '0',                  --      : IN  std_logic := '0';
--      s_axi_awready             =>  S_AXI_AWREADY,        --      : OUT std_logic;
--      s_axi_wid                 =>  "0000",         --(others => '0'),      --      : IN  std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_wdata               =>  "0000000000000000000000000000000000000000000000000000000000000000", --(others => '0'),      --      : IN  std_logic_vector(C_AXI_DATA_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_wstrb               =>  "00000000",          --(others => '0'),      --      : IN  std_logic_vector(C_AXI_DATA_WIDTH/8-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_wlast               =>  '0',                  --      : IN  std_logic := '0';
--      s_axi_wuser               =>  "0",            --(others => '0'),      --      : IN  std_logic_vector(C_AXI_WUSER_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_wvalid              =>  '0',                  --      : IN  std_logic := '0';
--      s_axi_wready              =>  S_AXI_WREADY,         --      : OUT std_logic;
--      s_axi_bid                 =>  S_AXI_BID,            --      : OUT std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_bresp               =>  S_AXI_BRESP,          --      : OUT std_logic_vector(2-1 DOWNTO 0);
--      s_axi_buser               =>  S_AXI_BUSER,          --      : OUT std_logic_vector(C_AXI_BUSER_WIDTH-1 DOWNTO 0);
--      s_axi_bvalid              =>  S_AXI_BVALID,          --      : OUT std_logic;
--      s_axi_bready              =>  '0',                  --      : IN  std_logic := '0';
--
--      -- AXI Full/Lite Master Write Channel (Read side)
--      m_axi_awid                =>  M_AXI_AWID,           --       : OUT std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0);
--      m_axi_awaddr              =>  M_AXI_AWADDR,         --       : OUT std_logic_vector(C_AXI_ADDR_WIDTH-1 DOWNTO 0);
--      m_axi_awlen               =>  M_AXI_AWLEN,          --       : OUT std_logic_vector(8-1 DOWNTO 0);
--      m_axi_awsize              =>  M_AXI_AWSIZE,         --       : OUT std_logic_vector(3-1 DOWNTO 0);
--      m_axi_awburst             =>  M_AXI_AWBURST,        --       : OUT std_logic_vector(2-1 DOWNTO 0);
--      m_axi_awlock              =>  M_AXI_AWLOCK,         --       : OUT std_logic_vector(2-1 DOWNTO 0);
--      m_axi_awcache             =>  M_AXI_AWCACHE,        --       : OUT std_logic_vector(4-1 DOWNTO 0);
--      m_axi_awprot              =>  M_AXI_AWPROT,         --       : OUT std_logic_vector(3-1 DOWNTO 0);
--      m_axi_awqos               =>  M_AXI_AWQOS,          --       : OUT std_logic_vector(4-1 DOWNTO 0);
--      m_axi_awregion            =>  M_AXI_AWREGION,       --       : OUT std_logic_vector(4-1 DOWNTO 0);
--      m_axi_awuser              =>  M_AXI_AWUSER,         --       : OUT std_logic_vector(C_AXI_AWUSER_WIDTH-1 DOWNTO 0);
--      m_axi_awvalid             =>  M_AXI_AWVALID,        --       : OUT std_logic;
--      m_axi_awready             =>  '0',                  --       : IN  std_logic := '0';
--      m_axi_wid                 =>  M_AXI_WID,            --       : OUT std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0);
--      m_axi_wdata               =>  M_AXI_WDATA,          --       : OUT std_logic_vector(C_AXI_DATA_WIDTH-1 DOWNTO 0);
--      m_axi_wstrb               =>  M_AXI_WSTRB,          --       : OUT std_logic_vector(C_AXI_DATA_WIDTH/8-1 DOWNTO 0);
--      m_axi_wlast               =>  M_AXI_WLAST,          --       : OUT std_logic;
--      m_axi_wuser               =>  M_AXI_WUSER,          --       : OUT std_logic_vector(C_AXI_WUSER_WIDTH-1 DOWNTO 0);
--      m_axi_wvalid              =>  M_AXI_WVALID,         --       : OUT std_logic;
--      m_axi_wready              =>  '0',                  --       : IN  std_logic := '0';
--      m_axi_bid                 =>  "0000",               --(others => '0'),      --       : IN  std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      m_axi_bresp               =>  "00",                 --(others => '0'),      --       : IN  std_logic_vector(2-1 DOWNTO 0) := (OTHERS => '0');
--      m_axi_buser               =>  "0",                  --(others => '0'),      --       : IN  std_logic_vector(C_AXI_BUSER_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      m_axi_bvalid              =>  '0',                  --       : IN  std_logic := '0';
--      m_axi_bready              =>  M_AXI_BREADY,         --       : OUT std_logic;
--
--      -- AXI Full/Lite Slave Read Channel (Write side)
--      s_axi_arid               =>  "0000",         --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_araddr             =>  "00000000000000000000000000000000",   --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(C_AXI_ADDR_WIDTH-1 DOWNTO 0) := (OTHERS => '0'); 
--      s_axi_arlen              =>  "00000000",          --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(8-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_arsize             =>  "000",          --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(3-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_arburst            =>  "00",           --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(2-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_arlock             =>  "00",           --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(2-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_arcache            =>  "0000",         --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(4-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_arprot             =>  "000",          --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(3-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_arqos              =>  "0000",         --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(4-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_arregion           =>  "0000",         --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(4-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_aruser             =>  "0",            --(others => '0'),      (others => '0'),       --       : IN  std_logic_vector(C_AXI_ARUSER_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axi_arvalid            =>  '0',                   --       : IN  std_logic := '0';
--      s_axi_arready            =>  S_AXI_ARREADY,         --       : OUT std_logic;
--      s_axi_rid                =>  S_AXI_RID,             --       : OUT std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0);       
--      s_axi_rdata              =>  S_AXI_RDATA,           --       : OUT std_logic_vector(C_AXI_DATA_WIDTH-1 DOWNTO 0); 
--      s_axi_rresp              =>  S_AXI_RRESP,           --       : OUT std_logic_vector(2-1 DOWNTO 0);
--      s_axi_rlast              =>  S_AXI_RLAST,           --       : OUT std_logic;
--      s_axi_ruser              =>  S_AXI_RUSER,           --       : OUT std_logic_vector(C_AXI_RUSER_WIDTH-1 DOWNTO 0);
--      s_axi_rvalid             =>  S_AXI_RVALID,          --       : OUT std_logic;
--      s_axi_rready             =>  '0',                   --       : IN  std_logic := '0';
--
--      -- AXI Full/Lite Master Read Channel (Read side)
--      m_axi_arid               =>  M_AXI_ARID,           --        : OUT std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0);        
--      m_axi_araddr             =>  M_AXI_ARADDR,         --        : OUT std_logic_vector(C_AXI_ADDR_WIDTH-1 DOWNTO 0);  
--      m_axi_arlen              =>  M_AXI_ARLEN,          --        : OUT std_logic_vector(8-1 DOWNTO 0);
--      m_axi_arsize             =>  M_AXI_ARSIZE,         --        : OUT std_logic_vector(3-1 DOWNTO 0);
--      m_axi_arburst            =>  M_AXI_ARBURST,        --        : OUT std_logic_vector(2-1 DOWNTO 0);
--      m_axi_arlock             =>  M_AXI_ARLOCK,         --        : OUT std_logic_vector(2-1 DOWNTO 0);
--      m_axi_arcache            =>  M_AXI_ARCACHE,        --        : OUT std_logic_vector(4-1 DOWNTO 0);
--      m_axi_arprot             =>  M_AXI_ARPROT,         --        : OUT std_logic_vector(3-1 DOWNTO 0);
--      m_axi_arqos              =>  M_AXI_ARQOS,          --        : OUT std_logic_vector(4-1 DOWNTO 0);
--      m_axi_arregion           =>  M_AXI_ARREGION,       --        : OUT std_logic_vector(4-1 DOWNTO 0);
--      m_axi_aruser             =>  M_AXI_ARUSER,         --        : OUT std_logic_vector(C_AXI_ARUSER_WIDTH-1 DOWNTO 0);
--      m_axi_arvalid            =>  M_AXI_ARVALID,        --        : OUT std_logic;
--      m_axi_arready            =>  '0',                  --        : IN  std_logic := '0';
--      m_axi_rid                =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_AXI_ID_WIDTH-1 DOWNTO 0) := (OTHERS => '0');        
--      m_axi_rdata              =>  "0000000000000000000000000000000000000000000000000000000000000000", --(others => '0'),      --        : IN  std_logic_vector(C_AXI_DATA_WIDTH-1 DOWNTO 0) := (OTHERS => '0');  
--      m_axi_rresp              =>  "00",                 --(others => '0'),      --        : IN  std_logic_vector(2-1 DOWNTO 0) := (OTHERS => '0');
--      m_axi_rlast              =>  '0',                  --        : IN  std_logic := '0';
--      m_axi_ruser              =>  "0",                  --(others => '0'),      --        : IN  std_logic_vector(C_AXI_RUSER_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      m_axi_rvalid             =>  '0',                  --        : IN  std_logic := '0';
--      m_axi_rready             =>  M_AXI_RREADY,         --        : OUT std_logic;
--
--      -- AXI Streaming Slave Signals (Write side)
--      s_axis_tvalid            =>  '0',                  --        : IN  std_logic := '0';
--      s_axis_tready            =>  S_AXIS_TREADY,        --        : OUT std_logic;
--      s_axis_tdata             =>  "0000000000000000000000000000000000000000000000000000000000000000", --(others => '0'),      --        : IN  std_logic_vector(C_AXIS_TDATA_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axis_tstrb             =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_AXIS_TSTRB_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axis_tkeep             =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_AXIS_TKEEP_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axis_tlast             =>  '0',                  --        : IN  std_logic := '0';
--      s_axis_tid               =>  "00000000",                 --(others => '0'),      --        : IN  std_logic_vector(C_AXIS_TID_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axis_tdest             =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_AXIS_TDEST_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--      s_axis_tuser             =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_AXIS_TUSER_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
--
--      -- AXI Streaming Master Signals (Read side)
--      m_axis_tvalid            =>  M_AXIS_TVALID,        --        : OUT std_logic;
--      m_axis_tready            =>  '0',                  --        : IN  std_logic := '0';
--      m_axis_tdata             =>  M_AXIS_TDATA,         --        : OUT std_logic_vector(C_AXIS_TDATA_WIDTH-1 DOWNTO 0);
--      m_axis_tstrb             =>  M_AXIS_TSTRB,         --        : OUT std_logic_vector(C_AXIS_TSTRB_WIDTH-1 DOWNTO 0);
--      m_axis_tkeep             =>  M_AXIS_TKEEP,         --        : OUT std_logic_vector(C_AXIS_TKEEP_WIDTH-1 DOWNTO 0);
--      m_axis_tlast             =>  M_AXIS_TLAST,         --        : OUT std_logic;
--      m_axis_tid               =>  M_AXIS_TID,           --        : OUT std_logic_vector(C_AXIS_TID_WIDTH-1 DOWNTO 0);
--      m_axis_tdest             =>  M_AXIS_TDEST,         --        : OUT std_logic_vector(C_AXIS_TDEST_WIDTH-1 DOWNTO 0);
--      m_axis_tuser             =>  M_AXIS_TUSER,         --        : OUT std_logic_vector(C_AXIS_TUSER_WIDTH-1 DOWNTO 0);
--
--      -- AXI Full/Lite Write Address Channel Signals
--      axi_aw_injectsbiterr     =>  '0',                  --        : IN  std_logic := '0';
--      axi_aw_injectdbiterr     =>  '0',                  --        : IN  std_logic := '0';
--      axi_aw_prog_full_thresh  =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_WR_PNTR_WIDTH_WACH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_aw_prog_empty_thresh =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_WR_PNTR_WIDTH_WACH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_aw_data_count        =>  AXI_AW_DATA_COUNT,    --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_WACH DOWNTO 0);
--      axi_aw_wr_data_count     =>  AXI_AW_WR_DATA_COUNT, --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_WACH DOWNTO 0);
--      axi_aw_rd_data_count     =>  AXI_AW_RD_DATA_COUNT, --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_WACH DOWNTO 0);
--      axi_aw_sbiterr           =>  AXI_AW_SBITERR,       --        : OUT std_logic;
--      axi_aw_dbiterr           =>  AXI_AW_DBITERR,       --        : OUT std_logic;
--      axi_aw_overflow          =>  AXI_AW_OVERFLOW,      --        : OUT std_logic;
--      axi_aw_underflow         =>  AXI_AW_UNDERFLOW,     --        : OUT std_logic;
--      axi_aw_prog_full         =>  AXI_AW_PROG_FULL,     --        : OUT STD_LOGIC := '0';
--      axi_aw_prog_empty        =>  AXI_AW_PROG_EMPTY,    --        : OUT STD_LOGIC := '1';
--
--
--      -- AXI Full/Lite Write Data Channel Signals
--      axi_w_injectsbiterr      =>  '0',                  --        : IN  std_logic := '0';
--      axi_w_injectdbiterr      =>  '0',                  --        : IN  std_logic := '0';
--      axi_w_prog_full_thresh   =>  "0000000000",         --(others => '0'),      --        : IN  std_logic_vector(C_WR_PNTR_WIDTH_WDCH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_w_prog_empty_thresh  =>  "0000000000",         --(others => '0'),      --        : IN  std_logic_vector(C_WR_PNTR_WIDTH_WDCH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_w_data_count         =>  AXI_W_DATA_COUNT,     --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_WDCH DOWNTO 0);
--      axi_w_wr_data_count      =>  AXI_W_WR_DATA_COUNT,  --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_WDCH DOWNTO 0);
--      axi_w_rd_data_count      =>  AXI_W_RD_DATA_COUNT,  --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_WDCH DOWNTO 0);
--      axi_w_sbiterr            =>  AXI_W_SBITERR,        --        : OUT std_logic;
--      axi_w_dbiterr            =>  AXI_W_DBITERR,        --        : OUT std_logic;
--      axi_w_overflow           =>  AXI_W_OVERFLOW,       --        : OUT std_logic;
--      axi_w_underflow          =>  AXI_W_UNDERFLOW,      --        : OUT std_logic;
--      axi_w_prog_full          =>  AXI_W_PROG_FULL,      --        : OUT STD_LOGIC := '0';
--      axi_w_prog_empty         =>  AXI_W_PROG_EMPTY,     --        : OUT STD_LOGIC := '1';
--
--      -- AXI Full/Lite Write Response Channel Signals
--      axi_b_injectsbiterr      =>  '0',                  --        : IN  std_logic := '0';
--      axi_b_injectdbiterr      =>  '0',                  --        : IN  std_logic := '0';
--      axi_b_prog_full_thresh   =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_WR_PNTR_WIDTH_WRCH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_b_prog_empty_thresh  =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_WR_PNTR_WIDTH_WRCH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_b_data_count         =>  AXI_B_DATA_COUNT,     --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_WRCH DOWNTO 0);
--      axi_b_wr_data_count      =>  AXI_B_WR_DATA_COUNT,  --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_WRCH DOWNTO 0);
--      axi_b_rd_data_count      =>  AXI_B_RD_DATA_COUNT,  --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_WRCH DOWNTO 0);
--      axi_b_sbiterr            =>  AXI_B_SBITERR,        --        : OUT std_logic;
--      axi_b_dbiterr            =>  AXI_B_DBITERR,        --        : OUT std_logic;
--      axi_b_overflow           =>  AXI_B_OVERFLOW,       --        : OUT std_logic;
--      axi_b_underflow          =>  AXI_B_UNDERFLOW,      --        : OUT std_logic;
--      axi_b_prog_full          =>  AXI_B_PROG_FULL,      --        : OUT STD_LOGIC := '0';
--      axi_b_prog_empty         =>  AXI_B_PROG_EMPTY,     --        : OUT STD_LOGIC := '1';
--
--      -- AXI Full/Lite Read Address Channel Signals
--      axi_ar_injectsbiterr     =>  '0',                  --        : IN  std_logic := '0';
--      axi_ar_injectdbiterr     =>  '0',                  --        : IN  std_logic := '0';
--      axi_ar_prog_full_thresh  =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_WR_PNTR_WIDTH_RACH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_ar_prog_empty_thresh =>  "0000",               --(others => '0'),      --        : IN  std_logic_vector(C_WR_PNTR_WIDTH_RACH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_ar_data_count        =>  AXI_AR_DATA_COUNT,    --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_RACH DOWNTO 0);
--      axi_ar_wr_data_count     =>  AXI_AR_WR_DATA_COUNT, --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_RACH DOWNTO 0);
--      axi_ar_rd_data_count     =>  AXI_AR_RD_DATA_COUNT, --        : OUT std_logic_vector(C_WR_PNTR_WIDTH_RACH DOWNTO 0);
--      axi_ar_sbiterr           =>  AXI_AR_SBITERR,       --        : OUT std_logic;
--      axi_ar_dbiterr           =>  AXI_AR_DBITERR,       --        : OUT std_logic;
--      axi_ar_overflow          =>  AXI_AR_OVERFLOW,      --        : OUT std_logic;
--      axi_ar_underflow         =>  AXI_AR_UNDERFLOW,     --        : OUT std_logic;
--      axi_ar_prog_full         =>  AXI_AR_PROG_FULL,     --        : OUT STD_LOGIC := '0';
--      axi_ar_prog_empty        =>  AXI_AR_PROG_EMPTY,    --        : OUT STD_LOGIC := '1';
--
--      -- AXI Full/Lite Read Data Channel Signals
--      axi_r_injectsbiterr     =>  '0',                  --         : IN  std_logic := '0';
--      axi_r_injectdbiterr     =>  '0',                  --         : IN  std_logic := '0';
--      axi_r_prog_full_thresh  =>  "0000000000",         --(others => '0'),      --         : IN  std_logic_vector(C_WR_PNTR_WIDTH_RDCH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_r_prog_empty_thresh =>  "0000000000",         --(others => '0'),      --         : IN  std_logic_vector(C_WR_PNTR_WIDTH_RDCH-1 DOWNTO 0) := (OTHERS => '0');
--      axi_r_data_count        =>  AXI_R_DATA_COUNT,     --         : OUT std_logic_vector(C_WR_PNTR_WIDTH_RDCH DOWNTO 0);
--      axi_r_wr_data_count     =>  AXI_R_WR_DATA_COUNT,  --         : OUT std_logic_vector(C_WR_PNTR_WIDTH_RDCH DOWNTO 0);
--      axi_r_rd_data_count     =>  AXI_R_RD_DATA_COUNT,  --         : OUT std_logic_vector(C_WR_PNTR_WIDTH_RDCH DOWNTO 0);
--      axi_r_sbiterr           =>  AXI_R_SBITERR,        --         : OUT std_logic;
--      axi_r_dbiterr           =>  AXI_R_DBITERR,        --         : OUT std_logic;
--      axi_r_overflow          =>  AXI_R_OVERFLOW,       --         : OUT std_logic;
--      axi_r_underflow         =>  AXI_R_UNDERFLOW,      --         : OUT std_logic;
--      axi_r_prog_full         =>  AXI_R_PROG_FULL,      --         : OUT STD_LOGIC := '0';
--      axi_r_prog_empty        =>  AXI_R_PROG_EMPTY,     --         : OUT STD_LOGIC := '1';
--
--      -- AXI Streaming FIFO Related Signals
--      axis_injectsbiterr      =>  '0',                  --         : IN  std_logic := '0';
--      axis_injectdbiterr      =>  '0',                  --         : IN  std_logic := '0';
--      axis_prog_full_thresh   =>  "0000000000",         --(others => '0'),      --         : IN  std_logic_vector(C_WR_PNTR_WIDTH_AXIS-1 DOWNTO 0) := (OTHERS => '0');
--      axis_prog_empty_thresh  =>  "0000000000",         --(others => '0'),      --         : IN  std_logic_vector(C_WR_PNTR_WIDTH_AXIS-1 DOWNTO 0) := (OTHERS => '0');
--      axis_data_count         =>  AXIS_DATA_COUNT,      --         : OUT std_logic_vector(C_WR_PNTR_WIDTH_AXIS DOWNTO 0);
--      axis_wr_data_count      =>  AXIS_WR_DATA_COUNT,   --         : OUT std_logic_vector(C_WR_PNTR_WIDTH_AXIS DOWNTO 0);
--      axis_rd_data_count      =>  AXIS_RD_DATA_COUNT,   --         : OUT std_logic_vector(C_WR_PNTR_WIDTH_AXIS DOWNTO 0);
--      axis_sbiterr            =>  AXIS_SBITERR,         --         : OUT std_logic;
--      axis_dbiterr            =>  AXIS_DBITERR,         --         : OUT std_logic;
--      axis_overflow           =>  AXIS_OVERFLOW,        --         : OUT std_logic;
--      axis_underflow          =>  AXIS_UNDERFLOW,       --         : OUT std_logic
--      axis_prog_full          =>  AXIS_PROG_FULL,       --         : OUT STD_LOGIC := '0';
--      axis_prog_empty         =>  AXIS_PROG_EMPTY       --         : OUT STD_LOGIC := '1';
--
--
--     
--      );

      

end implementation;



------------------------------------------------------------------------
-- Title      : Package for the rx_if logic
-- Project    : Tri-Mode Ethernet FIFO
------------------------------------------------------------------------
-- File       : rx_if_pack.vhd
-- Author     : Xilinx Inc.
------------------------------------------------------------------------
-- (c) Copyright 2012 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
------------------------------------------------------------------------
-- Description:  This package contains all component declarations for
--               the entiries which make up the Rx I/F logic
------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;



package rx_if_pack is


  component rx_if
  generic (
    C_FAMILY              : string                        := "virtex6";
    C_HAS_SGMII           : integer range 0 to 1          := 0;
    C_RXCSUM              : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_RXMEM               : integer                       := 4096;
    C_RXVLAN_TRAN         : integer range 0 to 1          := 0;
    C_RXVLAN_TAG          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP         : integer range 0 to 1          := 0;
    C_ENABLE_1588         : integer   := 0;
    C_MCAST_EXTEND        : integer range 0 to 1          := 0
    );

  port    (
    RX_FRAME_RECEIVED_INTRPT        : out std_logic;                          --  Frame received interrupt
    RX_FRAME_REJECTED_INTRPT        : out std_logic;                          --  Frame rejected interrupt
    RX_BUFFER_MEM_OVERFLOW_INTRPT   : out std_logic;                          --  Memory overflow interrupt

    AXI_STR_RXD_ACLK                : in  std_logic;                          --  AXI-Stream Receive Data Clock
    AXI_STR_RXD_VALID               : out std_logic;                          --  AXI-Stream Receive Data Valid
    AXI_STR_RXD_READY               : in  std_logic;                          --  AXI-Stream Receive Data Ready
    AXI_STR_RXD_LAST                : out std_logic;                          --  AXI-Stream Receive Data Last
    AXI_STR_RXD_STRB                : out std_logic_vector(3 downto 0);       --  AXI-Stream Receive Data Keep
    AXI_STR_RXD_DATA                : out std_logic_vector(31 downto 0);      --  AXI-Stream Receive Data Data
    RESET2AXI_STR_RXD               : in  std_logic;                          --  AXI-Stream Receive Data Reset

    AXI_STR_RXS_ACLK                : in  std_logic;                          --  AXI-Stream Receive Status Clock
    AXI_STR_RXS_VALID               : out std_logic;                          --  AXI-Stream Receive Status Valid
    AXI_STR_RXS_READY               : in  std_logic;                          --  AXI-Stream Receive Status Ready
    AXI_STR_RXS_LAST                : out std_logic;                          --  AXI-Stream Receive Status Last
    AXI_STR_RXS_STRB                : out std_logic_vector(3 downto 0);       --  AXI-Stream Receive Status Keep
    AXI_STR_RXS_DATA                : out std_logic_vector(31 downto 0);      --  AXI-Stream Receive Status Data
    RESET2AXI_STR_RXS               : in  std_logic;                          --  AXI-Stream Receive Status Reset

    -- added 05/5/2011
    RX_CLK_ENABLE_IN                : in std_logic;                           -- TEMAC clock domain enable

    rx_statistics_vector            : in  std_logic_vector(27 downto 0);      -- RX statistics from TEMAC
    rx_statistics_valid             : in  std_logic;                          -- Rx stats valid from TEMAC
    rxspeedis10100                  : in  std_logic;                          -- speed is 10/100 not 1000 indicator

    rx_mac_aclk                     : in  std_logic;                          -- Rx axistream clock from TEMAC
    rx_reset                        : in  std_logic;                          -- Rx axistream reset from TEMAC
    rx_axis_mac_tdata               : in  std_logic_vector(7 downto 0);       -- Rx axistream data from TEMAC
    rx_axis_mac_tvalid              : in  std_logic;                          -- Rx axistream valid from TEMAC
    rx_axis_mac_tlast               : in  std_logic;                          -- Rx axistream last from TEMAC
    rx_axis_mac_tuser               : in  std_logic;                          -- Rx axistream good/bad indicator from TEMAC

    RX_CL_CLK_RX_TAG_REG_DATA       : in  std_logic_vector(0 to 31);          --  Receive VLAN TAG
    RX_CL_CLK_TPID0_REG_DATA        : in  std_logic_vector(0 to 31);          --  Receive VLAN TPID 0
    RX_CL_CLK_TPID1_REG_DATA        : in  std_logic_vector(0 to 31);          --  Receive VLAN TPID 1
    RX_CL_CLK_UAWL_REG_DATA         : in  std_logic_vector(0 to 31);          --  Receive Unicast Address Word Lower
    RX_CL_CLK_UAWU_REG_DATA         : in  std_logic_vector(16 to 31);         --  Receive Unicast Address Word Upper

    RX_CL_CLK_MCAST_ADDR            : out std_logic_vector(0 to 14);          --  Receive Multicast Memory Address
    RX_CL_CLK_MCAST_EN              : out std_logic;                          --  Receive Multicast Memory Address Enable
    RX_CL_CLK_MCAST_RD_DATA         : in  std_logic_vector(0 to 0);           --  Receive Multicast Memory Address Read Data

    RX_CL_CLK_VLAN_ADDR             : out std_logic_vector(0 to 11);          --  Receive VLAN Memory Address
    RX_CL_CLK_VLAN_RD_DATA          : in  std_logic_vector(18 to 31);         --  Receive VLAN Memory Read Data
    RX_CL_CLK_VLAN_BRAM_EN_A        : out std_logic;                          --  Receive VLAN Memory Enable

    RX_CL_CLK_BAD_FRAME_ENBL        : in  std_logic;                          --  Receive Bad Frame Enable
    RX_CL_CLK_EMULTI_FLTR_ENBL      : in  std_logic;                          --  Receive Extended Multicast Address Filter Enable
    RX_CL_CLK_NEW_FNC_ENBL          : in  std_logic;                          --  Receive New Function Enable
    RX_CL_CLK_BRDCAST_REJ           : in  std_logic;                          --  Receive Broadcast Reject
    RX_CL_CLK_MULCAST_REJ           : in  std_logic;                          --  Receive Multicast Reject
    RX_CL_CLK_VSTRP_MODE            : in  std_logic_vector(0 to 1);           --  Receive VLAN Strip Mode
    RX_CL_CLK_VTAG_MODE             : in  std_logic_vector(0 to 1)            --  Receive VLAN TAG Mode

    );
  end component;


  component rx_emac_if_vlan
  generic (
    C_RXVLAN_WIDTH        : integer                       := 12;
    C_RXD_MEM_BYTES       : integer                       := 4096;
    C_RXD_MEM_ADDR_WIDTH  : integer                       := 10;
    C_RXS_MEM_BYTES       : integer                       := 4096;
    C_RXS_MEM_ADDR_WIDTH  : integer                       := 10;
    C_FAMILY              : string                        := "virtex6";
    C_RXCSUM              : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_RXVLAN_TRAN         : integer range 0 to 1          := 0;
    C_RXVLAN_TAG          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP         : integer range 0 to 1          := 0;
    C_MCAST_EXTEND        : integer range 0 to 1          := 0
    );

  port    (
    RX_FRAME_RECEIVED_INTRPT        : out std_logic;                        --  Frame received interrupt
    RX_FRAME_REJECTED_INTRPT        : out std_logic;                        --  Frame rejected interrupt
    RX_BUFFER_MEM_OVERFLOW_INTRPT   : out std_logic;                        --  Memory overflow interrupt

    rx_statistics_vector            : in  std_logic_vector(27 downto 0);
    rx_statistics_valid             : in  std_logic;
    end_of_frame_reset_in           : in  std_logic;

    rx_mac_aclk                     : in  std_logic;
    rx_reset                        : in  std_logic;
    derived_rxd                     : in  std_logic_vector(7 downto 0);

    derived_rx_good_frame           : in  std_logic;
    derived_rx_bad_frame            : in  std_logic;
    derived_rxd_vld                 : in  std_logic;
    derived_rx_clk_enbl             : in  std_logic;

    RX_CL_CLK_RX_TAG_REG_DATA       : in  std_logic_vector(0 to 31);        --  Receive VLAN TAG
    RX_CL_CLK_TPID0_REG_DATA        : in  std_logic_vector(0 to 31);        --  Receive VLAN TPID 0
    RX_CL_CLK_TPID1_REG_DATA        : in  std_logic_vector(0 to 31);        --  Receive VLAN TPID 1
    RX_CL_CLK_UAWL_REG_DATA         : in  std_logic_vector(0 to 31);        --  Receive Unicast Address Word Lower
    RX_CL_CLK_UAWU_REG_DATA         : in  std_logic_vector(16 to 31);       --  Receive Unicast Address Word Upper

    RX_CL_CLK_MCAST_ADDR            : out std_logic_vector(0 to 14);        --  Receive Multicast Memory Address
    RX_CL_CLK_MCAST_EN              : out std_logic;                        --  Receive Multicast Memory Address Enable
    RX_CL_CLK_MCAST_RD_DATA         : in  std_logic_vector(0 to 0);         --  Receive Multicast Memory Address Read Data

    RX_CL_CLK_VLAN_ADDR             : out std_logic_vector(0 to 11);        --  Receive VLAN Memory Address
    RX_CL_CLK_VLAN_RD_DATA          : in  std_logic_vector(18 to 31);       --  Receive VLAN Memory Read Data
    RX_CL_CLK_VLAN_BRAM_EN_A        : out std_logic;                        --  Receive VLAN Memory Enable

    RX_CL_CLK_BAD_FRAME_ENBL        : in  std_logic;                        --  Receive Bad Frame Enable
    RX_CL_CLK_EMULTI_FLTR_ENBL      : in  std_logic;                        --  Receive Extended Multicast Address Filter Enable
    RX_CL_CLK_NEW_FNC_ENBL          : in  std_logic;                        --  Receive New Function Enable
    RX_CL_CLK_BRDCAST_REJ           : in  std_logic;                        --  Receive Broadcast Reject
    RX_CL_CLK_MULCAST_REJ           : in  std_logic;                        --  Receive Multicast Reject
    RX_CL_CLK_VSTRP_MODE            : in  std_logic_vector(0 to 1);         --  Receive VLAN Strip Mode
    RX_CL_CLK_VTAG_MODE             : in  std_logic_vector(0 to 1);         --  Receive VLAN TAG Mode

    RX_CLIENT_RXD_DPMEM_WR_DATA     : out std_logic_vector(35 downto 0);                    --  Receive Data Memory Write Data
    RX_CLIENT_RXD_DPMEM_RD_DATA     : in  std_logic_vector(35 downto 0);                    --  Receive Data Memory Read Data
    RX_CLIENT_RXD_DPMEM_WR_EN       : out std_logic_vector(0 downto 0);                     --  Receive Data Memory Write Enable
    RX_CLIENT_RXD_DPMEM_ADDR        : out std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  Receive Data Memory Address
    RX_CLIENT_RXS_DPMEM_WR_DATA     : out std_logic_vector(35 downto 0);                    --  Receive Status Memory Write Data
    RX_CLIENT_RXS_DPMEM_RD_DATA     : in  std_logic_vector(35 downto 0);                    --  Receive Status Memory Read Data
    RX_CLIENT_RXS_DPMEM_WR_EN       : out std_logic_vector(0 downto 0);                     --  Receive Status Memory Write Enable
    RX_CLIENT_RXS_DPMEM_ADDR        : out std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  Receive Status Memory Address

    AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY : in std_logic_vector(35 downto 0);    --  Receive Status Gray code pointer
    AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY : in std_logic_vector(35 downto 0)     --  Receive Data Gray code pointer
  );
  end component;


  component rx_emac_if
  generic (
    C_RXVLAN_WIDTH        : integer                       := 12;
    C_RXD_MEM_BYTES       : integer                       := 4096;
    C_RXD_MEM_ADDR_WIDTH  : integer                       := 10;
    C_RXS_MEM_BYTES       : integer                       := 4096;
    C_RXS_MEM_ADDR_WIDTH  : integer                       := 10;
    C_FAMILY              : string                        := "virtex6";
    C_RXCSUM              : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_RXVLAN_TRAN         : integer range 0 to 1          := 0;
    C_RXVLAN_TAG          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP         : integer range 0 to 1          := 0;
    C_ENABLE_1588         : integer   := 0;
    C_MCAST_EXTEND        : integer range 0 to 1          := 0
    );

  port    (
    RX_FRAME_RECEIVED_INTRPT        : out std_logic;                        --  Frame received interrupt
    RX_FRAME_REJECTED_INTRPT        : out std_logic;                        --  Frame rejected interrupt
    RX_BUFFER_MEM_OVERFLOW_INTRPT   : out std_logic;                        --  Memory overflow interrupt

    rx_statistics_vector            : in  std_logic_vector(27 downto 0);    -- RX statistics from TEMAC
    rx_statistics_valid             : in  std_logic;                        -- Rx stats valid from TEMAC
    end_of_frame_reset_in           : in  std_logic;                        -- end of frame reset base on last from rx axistream

    rx_mac_aclk                     : in  std_logic;                        -- Rx axistream clock from TEMAC
    rx_reset                        : in  std_logic;                        -- Rx axistream reset from TEMAC
    derived_rxd                     : in  std_logic_vector(7 downto 0);     -- Rx axistream data from TEMAC

    derived_rx_good_frame           : in  std_logic;                        -- derived good indicator
    derived_rx_bad_frame            : in  std_logic;                        -- derived bad indicator
    derived_rxd_vld                 : in  std_logic;                        -- derived data valid indicator
    derived_rx_clk_enbl             : in  std_logic;                        -- TEMAC clock domain enable

    RX_CL_CLK_RX_TAG_REG_DATA       : in  std_logic_vector(0 to 31);        --  Receive VLAN TAG
    RX_CL_CLK_TPID0_REG_DATA        : in  std_logic_vector(0 to 31);        --  Receive VLAN TPID 0
    RX_CL_CLK_TPID1_REG_DATA        : in  std_logic_vector(0 to 31);        --  Receive VLAN TPID 1
    RX_CL_CLK_UAWL_REG_DATA         : in  std_logic_vector(0 to 31);        --  Receive Unicast Address Word Lower
    RX_CL_CLK_UAWU_REG_DATA         : in  std_logic_vector(16 to 31);       --  Receive Unicast Address Word Upper

    RX_CL_CLK_MCAST_ADDR            : out std_logic_vector(0 to 14);        --  Receive Multicast Memory Address
    RX_CL_CLK_MCAST_EN              : out std_logic;                        --  Receive Multicast Memory Address Enable
    RX_CL_CLK_MCAST_RD_DATA         : in  std_logic_vector(0 to 0);         --  Receive Multicast Memory Address Read Data

    RX_CL_CLK_VLAN_ADDR             : out std_logic_vector(0 to 11);        --  Receive VLAN Memory Address
    RX_CL_CLK_VLAN_RD_DATA          : in  std_logic_vector(18 to 31);       --  Receive VLAN Memory Read Data
    RX_CL_CLK_VLAN_BRAM_EN_A        : out std_logic;                        --  Receive VLAN Memory Enable

    RX_CL_CLK_BAD_FRAME_ENBL        : in  std_logic;                        --  Receive Bad Frame Enable
    RX_CL_CLK_EMULTI_FLTR_ENBL      : in  std_logic;                        --  Receive Extended Multicast Address Filter Enable
    RX_CL_CLK_NEW_FNC_ENBL          : in  std_logic;                        --  Receive New Function Enable
    RX_CL_CLK_BRDCAST_REJ           : in  std_logic;                        --  Receive Broadcast Reject
    RX_CL_CLK_MULCAST_REJ           : in  std_logic;                        --  Receive Multicast Reject
    RX_CL_CLK_VSTRP_MODE            : in  std_logic_vector(0 to 1);         --  Receive VLAN Strip Mode
    RX_CL_CLK_VTAG_MODE             : in  std_logic_vector(0 to 1);         --  Receive VLAN TAG Mode

    RX_CLIENT_RXD_DPMEM_WR_DATA     : out std_logic_vector(35 downto 0);                    --  Receive Data Memory Write Data
    RX_CLIENT_RXD_DPMEM_RD_DATA     : in  std_logic_vector(35 downto 0);                    --  Receive Data Memory Read Data
    RX_CLIENT_RXD_DPMEM_WR_EN       : out std_logic_vector(0 downto 0);                     --  Receive Data Memory Write Enable
    RX_CLIENT_RXD_DPMEM_ADDR        : out std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  Receive Data Memory Address
    RX_CLIENT_RXS_DPMEM_WR_DATA     : out std_logic_vector(35 downto 0);                    --  Receive Status Memory Write Data
    RX_CLIENT_RXS_DPMEM_RD_DATA     : in  std_logic_vector(35 downto 0);                    --  Receive Status Memory Read Data
    RX_CLIENT_RXS_DPMEM_WR_EN       : out std_logic_vector(0 downto 0);                     --  Receive Status Memory Write Enable
    RX_CLIENT_RXS_DPMEM_ADDR        : out std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  Receive Status Memory Address

    AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY : in std_logic_vector(35 downto 0);    --  Receive Status Gray code pointer
    AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY : in std_logic_vector(35 downto 0)     --  Receive Data Gray code pointer
  );
  end component;


  component rx_csum_if
  port (
    CLK       : in  std_logic;
    CLK_ENBL  : in  std_logic;
    RST       : in  std_logic;
    INTRFRMRST: in  std_logic;
    CALC_ENBL : in  std_logic;
    WORD_ENBL : in  std_logic;
    DATA_IN   : in  std_logic_vector(15 downto 0);
    CSUM_VLD  : out std_logic;
    CSUM      : out std_logic_vector(15 downto 0)
    );
  end component;


  component rx_axistream_if
  generic (
    C_RXD_MEM_BYTES       : integer                       := 4096;
    C_RXD_MEM_ADDR_WIDTH  : integer                       := 10;
    C_RXS_MEM_BYTES       : integer                       := 4096;
    C_RXS_MEM_ADDR_WIDTH  : integer                       := 10;
    C_FAMILY              : string                        := "virtex6";
    C_RXCSUM              : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_RXVLAN_TRAN         : integer range 0 to 1          := 0;
    C_RXVLAN_TAG          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP         : integer range 0 to 1          := 0;
    C_MCAST_EXTEND        : integer range 0 to 1          := 0
    );

  port    (
    AXI_STR_RXD_ACLK                : in  std_logic;                                        --  Receive AXI-Stream Data Clock
    AXI_STR_RXD_VALID               : out std_logic;                                        --  Receive AXI-Stream Data VALID
    AXI_STR_RXD_READY               : in  std_logic;                                        --  Receive AXI-Stream Data READY
    AXI_STR_RXD_LAST                : out std_logic;                                        --  Receive AXI-Stream Data LAST
    AXI_STR_RXD_STRB                : out std_logic_vector(3 downto 0);                     --  Receive AXI-Stream Data STRB
    AXI_STR_RXD_DATA                : out std_logic_vector(31 downto 0);                    --  Receive AXI-Stream Data DATA
    RESET2AXI_STR_RXD               : in  std_logic;                                        --  Reset

    AXI_STR_RXS_ACLK                : in  std_logic;                                        --  Receive AXI-Stream Status Clock
    AXI_STR_RXS_VALID               : out std_logic;                                        --  Receive AXI-Stream Status VALID
    AXI_STR_RXS_READY               : in  std_logic;                                        --  Receive AXI-Stream Status READY
    AXI_STR_RXS_LAST                : out std_logic;                                        --  Receive AXI-Stream Status LAST
    AXI_STR_RXS_STRB                : out std_logic_vector(3 downto 0);                     --  Receive AXI-Stream Status STRB
    AXI_STR_RXS_DATA                : out std_logic_vector(31 downto 0);                    --  Receive AXI-Stream Status DATA
    RESET2AXI_STR_RXS               : in  std_logic;                                        --  Reset

    AXI_STR_RXD_DPMEM_WR_DATA       : out std_logic_vector(35 downto 0);                    --  Receive Data Memory Wr Data
    AXI_STR_RXD_DPMEM_RD_DATA       : in  std_logic_vector(35 downto 0);                    --  Receive Data Memory Rd Data
    AXI_STR_RXD_DPMEM_WR_EN         : out std_logic_vector(0 downto 0);                     --  Receive Data Memory Wr Enable
    AXI_STR_RXD_DPMEM_ADDR          : out std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  Receive Data Memory Addr

    AXI_STR_RXS_DPMEM_WR_DATA       : out std_logic_vector(35 downto 0);                    --  Receive Status Memory Wr Data
    AXI_STR_RXS_DPMEM_RD_DATA       : in  std_logic_vector(35 downto 0);                    --  Receive Status Memory Rd Data
    AXI_STR_RXS_DPMEM_WR_EN         : out std_logic_vector(0 downto 0);                     --  Receive Status Memory Wr Enable
    AXI_STR_RXS_DPMEM_ADDR          : out std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  Receive Status Memory Addr

    AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY : out std_logic_vector(35 downto 0);             --  Receive Status GRAY Pointer
    AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY : out std_logic_vector(35 downto 0)              --  Receive Data GRAY Pointer
    );
  end component;


  component rx_mem_if
  generic (
    C_RXD_MEM_BYTES      : integer    := 4096;
    C_RXD_MEM_ADDR_WIDTH : integer    := 10;
    C_RXS_MEM_BYTES      : integer    := 4096;
    C_RXS_MEM_ADDR_WIDTH : integer    := 10;
    C_FAMILY             : string     := "virtex6"
  );

  port    (
    AXI_STR_RXD_ACLK            : in  std_logic;                                        --  AXI-Stream Receive Data Clock
    AXI_STR_RXD_DPMEM_WR_DATA   : in  std_logic_vector(35 downto 0);                    --  AXI-Stream Receive Data Write Data
    AXI_STR_RXD_DPMEM_RD_DATA   : out std_logic_vector(35 downto 0);                    --  AXI-Stream Receive Data Read Data
    AXI_STR_RXD_DPMEM_WR_EN     : in  std_logic_vector(0 downto 0);                     --  AXI-Stream Receive Data Write Enable
    AXI_STR_RXD_DPMEM_ADDR      : in  std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  AXI-Stream Receive Data Address
    RESET2AXI_STR_RXD           : in  std_logic;                                        --  AXI-Stream Receive Data Rese

    AXI_STR_RXS_ACLK            : in  std_logic;                                        --  AXI-Stream Receive Status Clock
    AXI_STR_RXS_DPMEM_WR_DATA   : in  std_logic_vector(35 downto 0);                    --  AXI-Stream Receive Status Write Data
    AXI_STR_RXS_DPMEM_RD_DATA   : out std_logic_vector(35 downto 0);                    --  AXI-Stream Receive Status Read Data
    AXI_STR_RXS_DPMEM_WR_EN     : in  std_logic_vector(0 downto 0);                     --  AXI-Stream Receive Status Write Enable
    AXI_STR_RXS_DPMEM_ADDR      : in  std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  AXI-Stream Receive Status Address
    RESET2AXI_STR_RXS           : in  std_logic;                                        --  AXI-Stream Receive Status Rese

    RX_CLIENT_CLK               : in  std_logic;                                        --  Receive MAC Clock
    RX_CLIENT_CLK_ENBL          : in  std_logic;                                        --  Receive MAC Clock Enable
    RX_CLIENT_RXD_DPMEM_WR_DATA : in  std_logic_vector(35 downto 0);                    --  Receive MAC Data Memory Write Data
    RX_CLIENT_RXD_DPMEM_RD_DATA : out std_logic_vector(35 downto 0);                    --  Receive MAC Data Memory Read Data
    RX_CLIENT_RXD_DPMEM_WR_EN   : in  std_logic_vector(0 downto 0);                     --  Receive MAC Data Memory Write Enable
    RX_CLIENT_RXD_DPMEM_ADDR    : in  std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  Receive MAC Data Memory Address

    RX_CLIENT_RXS_DPMEM_WR_DATA : in  std_logic_vector(35 downto 0);                    --  Receive MAC Status Memory Write Data
    RX_CLIENT_RXS_DPMEM_RD_DATA : out std_logic_vector(35 downto 0);                    --  Receive MAC Status Memory Read Data
    RX_CLIENT_RXS_DPMEM_WR_EN   : in  std_logic_vector(0 downto 0);                     --  Receive MAC Status Memory Write Enable
    RX_CLIENT_RXS_DPMEM_ADDR    : in  std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  Receive MAC Status Memory Address
    RESET2RX_CLIENT         : in  std_logic                                             --  Receive MAC Reset
  );
  end component;


end rx_if_pack;


------------------------------------------------------------------------------
-- rx_csum_if.vhd
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--
------------------------------------------------------------------------------
-- Filename:        rx_csum_if.vhd
-- Version:         v2.00a
-- Description:
--
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:      DRP
-- History:
--
--  <initials>      <date>
-- ^^^^^^
--      Description of changes. If multiple lines are needed to fully describe
--      the changes made to the design, these lines should align with each other.
-- ~~~~~~
--
--  <initials>      <date>
-- ^^^^^^
--      More changes
-- ~~~~~~
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of : out   std_logic; port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Libraries used;
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.rx_if_pack.all;

entity rx_csum_if is
  port (
    CLK       : in  std_logic;
    CLK_ENBL  : in  std_logic;
    RST       : in  std_logic;
    INTRFRMRST: in  std_logic;
    CALC_ENBL : in  std_logic;
    WORD_ENBL : in  std_logic;
    DATA_IN   : in  std_logic_vector(15 downto 0);
    CSUM_VLD  : out std_logic;
    CSUM      : out std_logic_vector(15 downto 0)
    );
end entity;

architecture beh of rx_csum_if is

  signal checksum            : unsigned(16 downto 0);
  signal calcEnable_d1       : std_logic;
  signal wordEnable_d1       : std_logic;
  signal endOfEnablePulse    : std_logic;
  signal endOfEnablePulse_d1 : std_logic;
  signal dataIn_d1           : std_logic_vector(15 downto 0);
  signal byteCount           : unsigned(2 downto 0);

  begin

    ---------------------------------------------------------------------------
    --
    ---------------------------------------------------------------------------
    process(CLK)
      begin
        if(rising_edge(CLK)) then
          if(RST='1' or INTRFRMRST='1') then
            dataIn_d1   <= (others => '0');
          else
            if(CLK_ENBL='1') then
              dataIn_d1   <= DATA_IN;
            end if;
          end if;
        end if;
    end process;

    process(CLK)
      begin
        if(rising_edge(CLK)) then
          if(RST='1' or INTRFRMRST='1') then
            endOfEnablePulse    <= '0';
            endOfEnablePulse_d1 <= '0';
            calcEnable_d1       <= '0';
            wordEnable_d1       <= '0';
          else
            if(CLK_ENBL='1') then
              wordEnable_d1       <= WORD_ENBL;
              calcEnable_d1       <= CALC_ENBL;
              endOfEnablePulse    <= not(CALC_ENBL) and calcEnable_d1;
              endOfEnablePulse_d1 <= endOfEnablePulse;
            end if;
          end if;
        end if;
    end process;

    ---------------------------------------------------------------------------
    -- this is where the checksum is calculated
    ---------------------------------------------------------------------------

    process(clk)
      begin
        if(rising_edge(clk)) then
          if(rst='1') then
            checksum    <= (others => '0');
            byteCount   <= (others => '0');
          else
            if(CLK_ENBL='1') then
              if(calcEnable_d1='1') then
                if (byteCount < X"7" and wordEnable_d1 = '1') then
                  byteCount <= byteCount + 1;
                end if;
                if (byteCount = x"7" and wordEnable_d1 = '1') then
                  if ((checksum + unsigned('0' & dataIn_d1)) > X"ffff") then
                    checksum <= checksum + unsigned('0' & dataIn_d1) - X"ffff";
                  else
                    checksum <= checksum + unsigned('0' & dataIn_d1);
                  end if;
                end if;
              else
                checksum   <= (others => '0');
                byteCount  <= (others => '0');
              end if;
            end if;
          end if;
        end if;
    end process;

    CSUM_VLD <= endOfEnablePulse_d1;

    process(CLK)
      begin
        if(rising_edge(CLK)) then
          if(RST='1' or INTRFRMRST='1') then
            CSUM  <= (others => '0');
          else
            if(CLK_ENBL='1') then
              if (checksum(15 downto 0) = X"0000") then
                CSUM  <= X"ffff";
              else
                CSUM  <= std_logic_vector(checksum(15 downto 0));
              end if;
            end if;
          end if;
        end if;
    end process;

end beh;


------------------------------------------------------------------------------
-- rx_emac_if_vlan.vhd
------------------------------------------------------------------------------
-- (c) Copyright 2004-2009 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, rtlLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-- ------------------------------------------------------------------------------
--
------------------------------------------------------------------------------
-- Filename:        rx_emac_if_vlan.vhd
-- Version:         v1.00a
-- Description:     Receive interface between AXIStream and Temac
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to rtlrove
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:          MSH
--
--  MSH     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of : out   std_logic; port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Libraries used;
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.rx_if_pack.all;

library work;
use work.clock_cross_pack.all;

-------------------------------------------------------------------------------
-- Definition of Generics :
-------------------------------------------------------------------------------
-- System generics
--  C_FAMILY              -- Xilinx FPGA Family
--  C_RXD_MEM_BYTES               -- Depth of RX memory in Bytes
--  C_RXCSUM
--     0  No checksum offloading
--     1  Partial (legacy) checksum offloading
--     2  Full checksum offloading
--  C_RXVLAN_TRAN         -- Enable RX enhanced VLAN translation
--  C_RXVLAN_TAG          -- Enable RX enhanced VLAN taging
--  C_RXVLAN_STRP         -- Enable RX enhanced VLAN striping
--  C_MCAST_EXTEND        -- Enable RX extended multicast address filtering

-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Definition of Ports :
-------------------------------------------------------------------------------
--    BUS2IP_CLK
--    BUS2IP_RESET
--
--    AXI_STR_RXD_ACLK
--    AXI_STR_RXD_ARESET
--    AXI_STR_RXD_VALID
--    AXI_STR_RXD_READY
--    AXI_STR_RXD_LAST
--    AXI_STR_RXD_STRB
--    AXI_STR_RXD_DATA
--
--    AXI_STR_RXS_ACLK
--    AXI_STR_RXS_ARESET
--    AXI_STR_RXS_VALID
--    AXI_STR_RXS_READY
--    AXI_STR_RXS_LAST
--    AXI_STR_RXS_STRB
--    AXI_STR_RXS_DATA
--
--    EMAC_CLIENT_RXD_LEGACY
--    EMAC_CLIENT_RXD_VLD_LEGACY
--    EMAC_CLIENT_RX_GOODFRAME_LEGACY
--    EMAC_CLIENT_RX_BADFRAME_LEGACY
--    EMAC_CLIENT_RX_FRAMEDROP
--    LEGACY_RX_FILTER_MATCH
--
--    RX_CLIENT_CLK
--    RX_CLIENT_CLK_ENBL
--
--    EMAC_CLIENT_RX_STATS
--    EMAC_CLIENT_RX_STATS_VLD
--    EMAC_CLIENT_RX_STATS_BYTE_VLD
--    EMAC_CLIENT_RXD_VLD_2STATS
--    rx_statistics_vector
--
--    RTAGREGDATA
--    TPID0REGDATA
--    TPID1REGDATA
--    RX_CL_CLK_UAWL_REG_DATA
--    RX_CL_CLK_UAWU_REG_DATA
--    RXCLCLKMCASTADDR
--    RXCLCLKMCASTEN
--    RXCLCLKMCASTRDDATA
--    LLINKCLKVLANADDR
--    LLINKCLKVLANRDDATA
--    LLINKCLKRXVLANBRAMENA
--
--    LLINKCLKEMULTIFLTRENBL
--    LLINKCLKNEWFNCENBL
--    LLINKCLKRXVSTRPMODE
--    LLINKCLKRXVTAGMODE
-------------------------------------------------------------------------------
----                  Entity Section
-------------------------------------------------------------------------------

entity rx_emac_if_vlan is
  generic (
    C_RXVLAN_WIDTH        : integer                       := 12;
    C_RXD_MEM_BYTES       : integer                       := 4096;
    C_RXD_MEM_ADDR_WIDTH  : integer                       := 10;
    C_RXS_MEM_BYTES       : integer                       := 4096;
    C_RXS_MEM_ADDR_WIDTH  : integer                       := 10;
                C_ENABLE_1588          : integer   := 0;
    C_FAMILY              : string                        := "virtex6";
    C_RXCSUM              : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_RXVLAN_TRAN         : integer range 0 to 1          := 0;
    C_RXVLAN_TAG          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP         : integer range 0 to 1          := 0;
    C_MCAST_EXTEND        : integer range 0 to 1          := 0
    );

  port    (
    RX_FRAME_RECEIVED_INTRPT        : out std_logic;                        --  Frame received interrupt
    RX_FRAME_REJECTED_INTRPT        : out std_logic;                        --  Frame rejected interrupt
    RX_BUFFER_MEM_OVERFLOW_INTRPT   : out std_logic;                        --  Memory overflow interrupt

    rx_statistics_vector            : in  std_logic_vector(27 downto 0);
    rx_statistics_valid             : in  std_logic;
    end_of_frame_reset_in           : in  std_logic;

    rx_mac_aclk                     : in  std_logic;
    rx_reset                        : in  std_logic;
    derived_rxd                     : in  std_logic_vector(7 downto 0);

    derived_rx_good_frame           : in  std_logic;
    derived_rx_bad_frame            : in  std_logic;
    derived_rxd_vld                 : in  std_logic;
    derived_rx_clk_enbl             : in  std_logic;

    RX_CL_CLK_RX_TAG_REG_DATA       : in  std_logic_vector(0 to 31);        --  Receive VLAN TAG
    RX_CL_CLK_TPID0_REG_DATA        : in  std_logic_vector(0 to 31);        --  Receive VLAN TPID 0
    RX_CL_CLK_TPID1_REG_DATA        : in  std_logic_vector(0 to 31);        --  Receive VLAN TPID 1
    RX_CL_CLK_UAWL_REG_DATA         : in  std_logic_vector(0 to 31);        --  Receive Unicast Address Word Lower
    RX_CL_CLK_UAWU_REG_DATA         : in  std_logic_vector(16 to 31);       --  Receive Unicast Address Word Upper

    RX_CL_CLK_MCAST_ADDR            : out std_logic_vector(0 to 14);        --  Receive Multicast Memory Address
    RX_CL_CLK_MCAST_EN              : out std_logic;                        --  Receive Multicast Memory Address Enable
    RX_CL_CLK_MCAST_RD_DATA         : in  std_logic_vector(0 to 0);         --  Receive Multicast Memory Address Read Data

    RX_CL_CLK_VLAN_ADDR             : out std_logic_vector(0 to 11);        --  Receive VLAN Memory Address
    RX_CL_CLK_VLAN_RD_DATA          : in  std_logic_vector(18 to 31);       --  Receive VLAN Memory Read Data
    RX_CL_CLK_VLAN_BRAM_EN_A        : out std_logic;                        --  Receive VLAN Memory Enable

    RX_CL_CLK_BAD_FRAME_ENBL        : in  std_logic;                        --  Receive Bad Frame Enable
    RX_CL_CLK_EMULTI_FLTR_ENBL      : in  std_logic;                        --  Receive Extended Multicast Address Filter Enable
    RX_CL_CLK_NEW_FNC_ENBL          : in  std_logic;                        --  Receive New Function Enable
    RX_CL_CLK_BRDCAST_REJ           : in  std_logic;                        --  Receive Broadcast Reject
    RX_CL_CLK_MULCAST_REJ           : in  std_logic;                        --  Receive Multicast Reject
    RX_CL_CLK_VSTRP_MODE            : in  std_logic_vector(0 to 1);         --  Receive VLAN Strip Mode
    RX_CL_CLK_VTAG_MODE             : in  std_logic_vector(0 to 1);         --  Receive VLAN TAG Mode

    RX_CLIENT_RXD_DPMEM_WR_DATA     : out std_logic_vector(35 downto 0);                    --  Receive Data Memory Write Data
    RX_CLIENT_RXD_DPMEM_RD_DATA     : in  std_logic_vector(35 downto 0);                    --  Receive Data Memory Read Data
    RX_CLIENT_RXD_DPMEM_WR_EN       : out std_logic_vector(0 downto 0);                     --  Receive Data Memory Write Enable
    RX_CLIENT_RXD_DPMEM_ADDR        : out std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  Receive Data Memory Address
    RX_CLIENT_RXS_DPMEM_WR_DATA     : out std_logic_vector(35 downto 0);                    --  Receive Status Memory Write Data
    RX_CLIENT_RXS_DPMEM_RD_DATA     : in  std_logic_vector(35 downto 0);                    --  Receive Status Memory Read Data
    RX_CLIENT_RXS_DPMEM_WR_EN       : out std_logic_vector(0 downto 0);                     --  Receive Status Memory Write Enable
    RX_CLIENT_RXS_DPMEM_ADDR        : out std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  Receive Status Memory Address

    AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY : in std_logic_vector(35 downto 0);    --  Receive Status Gray code pointer
    AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY : in std_logic_vector(35 downto 0)     --  Receive Data Gray code pointer
  );
end rx_emac_if_vlan;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of rx_emac_if_vlan is

signal EMAC_CLIENT_RXD_LEGACY          : std_logic_vector(7 downto  0);
signal EMAC_CLIENT_RXD_VLD_LEGACY      : std_logic;
signal EMAC_CLIENT_RX_GOODFRAME_LEGACY : std_logic;
signal EMAC_CLIENT_RX_BADFRAME_LEGACY  : std_logic;
signal EMAC_CLIENT_RX_FRAMEDROP        : std_logic;
signal LEGACY_RX_FILTER_MATCH          : std_logic_vector(7 downto 0);

signal RX_CLIENT_CLK                   : std_logic;
signal RX_CLIENT_CLK_ENBL              : std_logic;
signal RESET2RX_CLIENT                 : std_logic;

signal EMAC_CLIENT_RX_STATS            : std_logic_vector(6  downto  0);
signal EMAC_CLIENT_RX_STATS_VLD        : std_logic;
signal EMAC_CLIENT_RX_STATS_BYTE_VLD   : std_logic;
signal EMAC_CLIENT_RXD_VLD_2STATS      : std_logic;
signal SOFT_EMAC_CLIENT_RX_STATS       : std_logic_vector(27 downto 0);

---------------------------------------------------------------------
-- Functions
---------------------------------------------------------------------

-- Convert a gray code value into binary
function gray_to_bin (
   gray : std_logic_vector)
   return std_logic_vector is

   variable binary : std_logic_vector(gray'range);

begin

   for i in gray'high downto gray'low loop
      if i = gray'high then
         binary(i) := gray(i);
      else
         binary(i) := binary(i+1) xor gray(i);
      end if;
   end loop;  -- i

   return binary;

end gray_to_bin;

------------------------------------------------------------------------------
-- Constant Declarations
------------------------------------------------------------------------------


------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

type type_rx_data_words_array    is array (1 to 8) of std_logic_vector(31 downto 0);
type type_rx_data_valid_array    is array (1 to 8) of std_logic_vector(3 downto 0);
type type_rx_data_packed_ready   is array (1 to 8) of std_logic;
type type_start_of_frame_array   is array (1 to 29) of std_logic;
type type_end_of_frame_array     is array (1 to 5) of std_logic;
type type_rx_data_packed_ready_array is array (1 to 8) of std_logic;

type RECEIVE_FRAME_CTRL_TYPE is (
          RESET_INIT_MEM_PTR_1,
          RESET_INIT_MEM_PTR_2,
          RESET_INIT_MEM_PTR_3,
          RESET_INIT_MEM_PTR_4,
          IDLE,
          UPDATE_MEM_PTR_1,
          UPDATE_STATUS_FIFO_WORD_1,
          UPDATE_STATUS_FIFO_WORD_2,
          UPDATE_STATUS_FIFO_WORD_3,
          UPDATE_STATUS_FIFO_WORD_4,
          UPDATE_STATUS_FIFO_WORD_5,
          UPDATE_STATUS_FIFO_WORD_6,
          UPDATE_MEM_PTR_2
        );

type RECEIVE_FRAME_DATA_TYPE is (
          RESET,
          WAIT_FOR_START_OF_FRAME,
          RECEIVING_FRAME,
          END_OF_FRAME_CHECK_GOOD_BAD
        );

signal receive_frame_current_state : RECEIVE_FRAME_CTRL_TYPE;
signal receive_frame_next_state    : RECEIVE_FRAME_CTRL_TYPE;

signal receive_frame_data_current_state : RECEIVE_FRAME_DATA_TYPE;
signal receive_frame_data_next_state    : RECEIVE_FRAME_DATA_TYPE;

signal rx_data_words_array    : type_rx_data_words_array;
signal rx_data_valid_array    : type_rx_data_valid_array;
signal start_of_frame_array   : type_start_of_frame_array;
signal end_of_frame_array     : type_end_of_frame_array;
signal rx_data_packed_ready_array : type_rx_data_packed_ready_array;

signal start_of_frame_d1    : std_logic;
signal save_rx_goodframe    : std_logic;
signal save_rx_badframe     : std_logic;


signal frame_is_multicast_d10           : std_logic;
signal frame_is_ip_multicast_d4         : std_logic;
signal frame_is_broadcast_d10           : std_logic;
signal frame_is_vlan_8100_d15           : std_logic;
signal first_tag_is_vlan_TPID_0_d15     : std_logic;
signal first_tag_is_vlan_TPID_1_d15     : std_logic;
signal first_tag_is_vlan_TPID_2_d15     : std_logic;
signal first_tag_is_vlan_TPID_3_d15     : std_logic;
signal second_tag_is_vlan_TPID_0_d19    : std_logic;
signal second_tag_is_vlan_TPID_1_d19    : std_logic;
signal second_tag_is_vlan_TPID_2_d19    : std_logic;
signal second_tag_is_vlan_TPID_3_d19    : std_logic;
signal frame_has_valid_length_field_d22 : std_logic;
signal frame_has_type_0800_d22          : std_logic;
signal frame_is_snap_d30                : std_logic;



signal rx_data_packed_word              : std_logic_vector(31 downto 0);
signal rx_data_vld_packed_word          : std_logic_vector(3 downto 0);
signal rx_data_packed_state             : unsigned(1 downto 0);
signal rx_data_packed_ready             : std_logic;

signal frame_length_bytes               : unsigned(15 downto 0);
signal frame_length_bytes_lat           : unsigned(15 downto 0);

signal rxd_mem_next_available4write_ptr_cmb : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_next_available4write_ptr_reg : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_last_read_out_ptr_cmb        : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_last_read_out_ptr_reg        : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_next_available4write_ptr_cmb : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_next_available4write_ptr_reg : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);

signal rxd_mem_full_mask                : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_full_mask_minus_one      : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_empty_mask               : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_one_mask                 : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_two_mask                 : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_full_mask                : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_full_mask_minus_one      : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_empty_mask               : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_one_mask                 : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_two_mask                 : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_three_mask               : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_four_mask                : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);

signal zero_extend_rxd_mask36           : std_logic_vector(35 downto C_RXD_MEM_ADDR_WIDTH + 1);
signal zero_extend_rxs_mask36           : std_logic_vector(35 downto C_RXS_MEM_ADDR_WIDTH + 1);

signal rxs_status_word_1_cmb            : std_logic_vector(35 downto 0);
signal rxs_status_word_1_reg            : std_logic_vector(35 downto 0);
signal rxs_status_word_2                : std_logic_vector(35 downto 0);
signal rxs_status_word_3                : std_logic_vector(35 downto 0);
signal rxs_status_word_4                : std_logic_vector(35 downto 0);
signal rxs_status_word_5                : std_logic_vector(35 downto 0);
signal rxs_status_word_6_cmb            : std_logic_vector(35 downto 0);
signal rxs_status_word_6_reg            : std_logic_vector(35 downto 0);

signal rxd_addr_cntr_en                 : std_logic;
signal rxs_addr_cntr_en                 : std_logic;
signal rxd_mem_addr_cntr                : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_addr_cntr                : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxd_addr_cntr_load               : std_logic;
signal rxs_addr_cntr_load               : std_logic;
signal update_status_fifo               : std_logic;

signal multicast_addr_upper_d10         : std_logic_vector(15 downto 0);
signal multicast_addr_lower_d10         : std_logic_vector(31 downto 0);
signal bytes_12_and_13_d19              : std_logic_vector(15 downto 0);
signal bytes_14_and_15_d19              : std_logic_vector(15 downto 0);

signal receive_checksum_status          : std_logic_vector(2 downto 0);
signal raw_checksum                     : std_logic_vector(15 downto 0);

signal statistics_vector                : std_logic_vector(25 downto 0);
signal frame_drop                       : std_logic;
signal not_enough_rxs_memory            : std_logic;

signal rxCsum                           : std_logic_vector(15 downto 0);
signal rxCsumVld                        : std_logic;
signal first_vlan_tag_vid_d17           : std_logic_vector(11 downto 0);
signal second_vlan_tag_vid_d21          : std_logic_vector(11 downto 0);
signal first_vlan_tag_bram_value_d18    : std_logic_vector(18 to 31);
signal second_vlan_tag_bram_value_d22   : std_logic_vector(18 to 31);
signal wd4TPIDMatch_d15                 : std_logic;
signal wd5TPIDMatch_d19                 : std_logic;
signal word4TagEnabled_d18              : std_logic;
signal word5TagEnabled_d22              : std_logic;
signal word4StrpEnabled_d18             : std_logic;
signal word4TransEnabled_d18            : std_logic;
signal word5TransEnabled_d19            : std_logic;
signal autoInsertWord4VlanTag           : std_logic;
signal autoInsertWord5VlanTag           : std_logic;
signal translateWord4VlanVid            : std_logic;
signal translateWord5VlanVid            : std_logic;
signal stripWord4VlanTag                : std_logic;
signal saveAutoInsertWord4VlanTag       : std_logic;
signal saveAutoInsertWord5VlanTag       : std_logic;
signal saveStripWord4VlanTag            : std_logic;
signal rx_cl_clk_vlan_addr_reg          : std_logic_vector(0 to 11);


signal extendedMulticastReject  : std_logic;
signal saveExtendedMulticastReject : std_logic;

signal rxclclk_rxd_mem_last_read_out_ptr           : std_logic_vector(35 downto 0);
signal rxclclk_rxd_mem_last_read_out_ptr_d1        : std_logic_vector(35 downto 0);
signal sync_rxd_mem_last_read_out_ptr_gray_sync    : std_logic_vector(35 downto 0);

signal rxclclk_rxs_mem_last_read_out_ptr           : std_logic_vector(35 downto 0);
signal rxclclk_rxs_mem_last_read_out_ptr_d1        : std_logic_vector(35 downto 0);
signal sync_rxs_mem_last_read_out_ptr_gray_sync      : std_logic_vector(35 downto 0);

signal eof_reset : std_logic;

signal initial_index       : integer;
begin

  EMAC_CLIENT_RXD_VLD_LEGACY      <= derived_rxd_vld;
  RX_CLIENT_CLK_ENBL              <= derived_rx_clk_enbl;

  EMAC_CLIENT_RX_GOODFRAME_LEGACY <= derived_rx_good_frame;
  EMAC_CLIENT_RX_BADFRAME_LEGACY  <= derived_rx_bad_frame;
  EMAC_CLIENT_RX_STATS_VLD        <= rx_statistics_valid;
  SOFT_EMAC_CLIENT_RX_STATS       <= rx_statistics_vector;
  RX_CLIENT_CLK                   <= rx_mac_aclk;
  RESET2RX_CLIENT                 <= rx_reset;
  EMAC_CLIENT_RXD_LEGACY          <= derived_rxd;

  eof_reset <= end_of_frame_reset_in;

    ENABLE_ZERO_INIT_CNT: if(C_ENABLE_1588 = 0) generate
    begin 
	initial_index <= 0;
    end generate ENABLE_ZERO_INIT_CNT;

    ENABLE_EIGHT_INIT_CNT: if(C_ENABLE_1588 > 0) generate
    begin 
	initial_index <= 8;
    end generate ENABLE_EIGHT_INIT_CNT;
  -------------------------------------------------------------------------
  -- Synchronize gray encoded last processed pointer from AXIStream clock
  -- domain to the receive client clock domain.
  -------------------------------------------------------------------------
  SYNC_RXS_LAST_READ_GRAY_PROCESS: for i in 35 downto 0 generate
     SYNC_RXS_LAST_READ_GRAY: sync_block
     port map (
        clk       => RX_CLIENT_CLK,
        reset     => RESET2RX_CLIENT,
        data_in   => AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY(i),
        data_out  => sync_rxs_mem_last_read_out_ptr_gray_sync(i)
     );
  end generate;


  -------------------------------------------------------------------------
  -- Convert gray encoded last processed pointer back to binary encoded
  -------------------------------------------------------------------------
  rxclclk_rxs_mem_last_read_out_ptr <= gray_to_bin(sync_rxs_mem_last_read_out_ptr_gray_sync);

  -------------------------------------------------------------------------
  -- Register binary encoded last processed pointer from local link
  -- interface
  -------------------------------------------------------------------------
  RX_CL_CLK_REG_RXS_LAST_READ_PROCESS: process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        rxclclk_rxs_mem_last_read_out_ptr_d1  <= (others => '0');
      else
        rxclclk_rxs_mem_last_read_out_ptr_d1  <= rxclclk_rxs_mem_last_read_out_ptr;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- Synchronize gray encoded last processed pointer from AXIStream clock
  -- domain to the receive client clock domain.
  -------------------------------------------------------------------------
  SYNC_RXD_LAST_READ_GRAY_PROCESS: for i in 35 downto 0 generate
     SYNC_RXD_LAST_READ_GRAY: sync_block
     port map (
        clk       => RX_CLIENT_CLK,
        reset     => RESET2RX_CLIENT,
        data_in   => AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY(i),
        data_out  => sync_rxd_mem_last_read_out_ptr_gray_sync(i)
     );
  end generate;

  -------------------------------------------------------------------------
  -- Convert gray encoded last processed pointer back to binary encoded
  -------------------------------------------------------------------------
  rxclclk_rxd_mem_last_read_out_ptr <= gray_to_bin(sync_rxd_mem_last_read_out_ptr_gray_sync);

  -------------------------------------------------------------------------
  -- Register binary encoded last processed pointer from local link
  -- interface
  -------------------------------------------------------------------------
  RX_CL_CLK_REG_RXD_LAST_READ_PROCESS: process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        rxclclk_rxd_mem_last_read_out_ptr_d1  <= (others => '0');
      else
        rxclclk_rxd_mem_last_read_out_ptr_d1  <= rxclclk_rxd_mem_last_read_out_ptr;
      end if;
    end if;
  end process;

  -----------------------------------------------------------------------------

  receive_checksum_status     <= (others => '0');

  rxs_status_word_2               <= X"00000" & multicast_addr_upper_d10;
  rxs_status_word_3               <= X"0" & multicast_addr_lower_d10;
  rxs_status_word_4               <= X"0" & statistics_vector & receive_checksum_status & frame_is_broadcast_d10 &
                                          frame_is_ip_multicast_d4 & frame_is_multicast_d10;
  rxs_status_word_5               <= X"0" & bytes_12_and_13_d19 & raw_checksum;
  rxs_status_word_6_cmb(35 downto 16) <= X"0" & bytes_14_and_15_d19;

  wd4TPIDMatch_d15 <= first_tag_is_vlan_TPID_0_d15 or first_tag_is_vlan_TPID_1_d15 or first_tag_is_vlan_TPID_2_d15 or first_tag_is_vlan_TPID_3_d15;
  wd5TPIDMatch_d19 <= second_tag_is_vlan_TPID_0_d19 or second_tag_is_vlan_TPID_1_d19 or second_tag_is_vlan_TPID_2_d19 or second_tag_is_vlan_TPID_3_d19;

  -------------------------------------------------------------------------
  -- Force extra write to memory
  -------------------------------------------------------------------------
  word4TagEnabled_d18 <= '1' when RX_CL_CLK_NEW_FNC_ENBL = '1' and C_RXVLAN_TAG  = 1 and
                                   ((RX_CL_CLK_VTAG_MODE = "01") or
                                    (RX_CL_CLK_VTAG_MODE = "10" and (word4StrpEnabled_d18 = '0' and wd4TPIDMatch_d15 = '1')) or
                                    (RX_CL_CLK_VTAG_MODE = "11" and ((word4StrpEnabled_d18 = '0' and wd4TPIDMatch_d15 = '1' and first_vlan_tag_bram_value_d18(31) = '1')))) else
                         '0';

  -------------------------------------------------------------------------
  -- Force extra write to memory
  -------------------------------------------------------------------------
  word5TagEnabled_d22 <= '1' when RX_CL_CLK_NEW_FNC_ENBL = '1' and C_RXVLAN_TAG  = 1 and
                                   ((RX_CL_CLK_VTAG_MODE = "10" and (word4StrpEnabled_d18 = '1' and wd5TPIDMatch_d19 = '1')) or
                                    (RX_CL_CLK_VTAG_MODE = "11" and ((word4StrpEnabled_d18 = '1' and wd5TPIDMatch_d19 = '1' and second_vlan_tag_bram_value_d22(31) = '1')))) else
                         '0';

  -------------------------------------------------------------------------
  -- Block write to memory
  -------------------------------------------------------------------------
  word4StrpEnabled_d18 <= '1' when RX_CL_CLK_NEW_FNC_ENBL = '1' and C_RXVLAN_STRP = 1 and
                                    ((RX_CL_CLK_VSTRP_MODE = "01" and wd4TPIDMatch_d15 = '1') or
                                     (RX_CL_CLK_VSTRP_MODE = "11" and wd4TPIDMatch_d15 = '1' and first_vlan_tag_bram_value_d18(30) = '1')) else
                          '0';

  -------------------------------------------------------------------------
  -- Substitute dat for write to memory
  -------------------------------------------------------------------------
  word4TransEnabled_d18 <= '1' when RX_CL_CLK_NEW_FNC_ENBL = '1' and C_RXVLAN_TRAN = 1 and
                                     ((word4StrpEnabled_d18 = '0' and wd4TPIDMatch_d15 = '1')) else
                           '0';

  -------------------------------------------------------------------------
  -- Substitute dat for write to memory
  -------------------------------------------------------------------------
  word5TransEnabled_d19 <= '1' when RX_CL_CLK_NEW_FNC_ENBL = '1' and C_RXVLAN_TRAN = 1 and
                                     ((word4StrpEnabled_d18 = '1' and wd5TPIDMatch_d19 = '1')) else
                           '0';

  -------------------------------------------------------------------------
  -- Generate variable width address masks for checking memory pointers
  -------------------------------------------------------------------------
  RXD_GEN_MASK: for I in C_RXD_MEM_ADDR_WIDTH downto 0 generate
    rxd_mem_full_mask(I) <= '1';
    rxd_mem_empty_mask(I)  <= '0';
  end generate;

  rxd_mem_one_mask            <= rxd_mem_empty_mask + 1;
  rxd_mem_two_mask            <= rxd_mem_empty_mask + 2;
  rxd_mem_full_mask_minus_one <= rxd_mem_full_mask - 1;

  RXS_GEN_MASK: for I in C_RXS_MEM_ADDR_WIDTH downto 0 generate
    rxs_mem_full_mask(I) <= '1';
    rxs_mem_empty_mask(I)  <= '0';
  end generate;

  rxs_mem_one_mask            <= rxs_mem_empty_mask + 1;
  rxs_mem_two_mask            <= rxs_mem_empty_mask + 2;
  rxs_mem_three_mask          <= rxs_mem_empty_mask + 3;
  rxs_mem_four_mask           <= rxs_mem_empty_mask + 4;
  rxs_mem_full_mask_minus_one <= rxs_mem_full_mask - 1;

  zero_extend_rxd_mask36      <= (others => '0');
  zero_extend_rxs_mask36      <= (others => '0');

  -------------------------------------------------------------------------
  -- pack the 8 bit wide client receive data into 32 bit wide
  -------------------------------------------------------------------------

  RX_DATA_8_TO_32_PACK : process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        rx_data_packed_word      <= (others => '0');
        rx_data_vld_packed_word  <= (others => '0');
        rx_data_packed_state     <= (others => '0');
        rx_data_packed_ready     <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (EMAC_CLIENT_RXD_VLD_LEGACY = '1') then -- word full and ready to use
            if (rx_data_packed_state = "11") then
              rx_data_packed_state <= (others => '0');
              rx_data_packed_ready <= '1';
            else
              rx_data_packed_state <= rx_data_packed_state + 1;
              rx_data_packed_ready <= '0';
            end if;
            if (rx_data_packed_state = "00") then
              rx_data_vld_packed_word(3)        <= EMAC_CLIENT_RXD_VLD_LEGACY;
              rx_data_packed_word(31 downto 24) <= EMAC_CLIENT_RXD_LEGACY;
            elsif(rx_data_packed_state = "01") then
              rx_data_vld_packed_word(3 downto 2) <= EMAC_CLIENT_RXD_VLD_LEGACY & rx_data_vld_packed_word(3);
              rx_data_packed_word(31 downto 16)   <= EMAC_CLIENT_RXD_LEGACY & rx_data_packed_word(31 downto 24);
            elsif(rx_data_packed_state = "10") then
              rx_data_vld_packed_word(3 downto 1) <= EMAC_CLIENT_RXD_VLD_LEGACY & rx_data_vld_packed_word(3 downto 2);
              rx_data_packed_word(31 downto 8)    <= EMAC_CLIENT_RXD_LEGACY     & rx_data_packed_word(31 downto 16);
            elsif(rx_data_packed_state = "11") then
              rx_data_vld_packed_word(3 downto 0) <= EMAC_CLIENT_RXD_VLD_LEGACY & rx_data_vld_packed_word(3 downto 1);
              rx_data_packed_word(31 downto 0)    <= EMAC_CLIENT_RXD_LEGACY     & rx_data_packed_word(31 downto 8);
            end if;
          elsif (EMAC_CLIENT_RXD_VLD_LEGACY = '0' and rx_data_valid_array(1)(0) = '1') then
            if(rx_data_packed_state = "01") then
              rx_data_vld_packed_word(3 downto 0) <= "000" & rx_data_vld_packed_word(3);
              rx_data_packed_word(31 downto 0)    <= "000000000000000000000000" & rx_data_packed_word(31 downto 24);
              rx_data_packed_ready <= '1';
              rx_data_packed_state     <= (others => '0');
            elsif(rx_data_packed_state = "10") then
              rx_data_vld_packed_word(3 downto 0) <= "00" & rx_data_vld_packed_word(3 downto 2);
              rx_data_packed_word(31 downto 0)    <= "0000000000000000" & rx_data_packed_word(31 downto 16);
              rx_data_packed_ready <= '1';
              rx_data_packed_state     <= (others => '0');
            elsif(rx_data_packed_state = "11") then
              rx_data_vld_packed_word(3 downto 0) <= '0' & rx_data_vld_packed_word(3 downto 1);
              rx_data_packed_word(31 downto 0)    <= "00000000" & rx_data_packed_word(31 downto 8);
              rx_data_packed_ready <= '1';
              rx_data_packed_state     <= (others => '0');
            else
              rx_data_packed_word      <= (others => '0');
              rx_data_vld_packed_word  <= (others => '0');
              rx_data_packed_state     <= (others => '0');
              rx_data_packed_ready     <= '0';
            end if;
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- calculate the partial checksum or not
  -------------------------------------------------------------------------

  INCLUDE_RX_CSUM: if(C_RXCSUM = 1) generate
    signal emacClientRxdLegacy_d1    : std_logic_vector(7 downto 0);
    signal rxd16bits                 : std_logic_vector(15 downto 0);
    signal emacClientRxdVldLegacy_d1 : std_logic;
    signal emacClientRxdVldWord      : std_logic;
  begin
    process(RX_CLIENT_CLK)
      begin
        if(rising_edge(RX_CLIENT_CLK)) then
          if(RESET2RX_CLIENT='1') then
            emacClientRxdLegacy_d1   <= (others => '0');
            emacClientRxdVldWord<= '0';
          else
            if(RX_CLIENT_CLK_ENBL='1') then
              emacClientRxdLegacy_d1   <= EMAC_CLIENT_RXD_LEGACY;
              emacClientRxdVldLegacy_d1<= EMAC_CLIENT_RXD_VLD_LEGACY;
              if (EMAC_CLIENT_RXD_VLD_LEGACY = '1' or emacClientRxdVldLegacy_d1 = '1') then
                emacClientRxdVldWord <= NOT(emacClientRxdVldWord);
              else
                emacClientRxdVldWord<= '0';
              end if;
            end if;
          end if;
        end if;
    end process;

    rxd16bits <= emacClientRxdLegacy_d1 & EMAC_CLIENT_RXD_LEGACY when EMAC_CLIENT_RXD_VLD_LEGACY = '1' else
                 emacClientRxdLegacy_d1 & X"00";

    I_RX_CSUM : rx_csum_if
      port map(
        CLK       => RX_CLIENT_CLK,
        CLK_ENBL  => RX_CLIENT_CLK_ENBL,
        RST       => RESET2RX_CLIENT,
        INTRFRMRST=> eof_reset,
        CALC_ENBL => emacClientRxdVldLegacy_d1,
        WORD_ENBL => emacClientRxdVldWord,
        DATA_IN   => rxd16bits,
        CSUM_VLD  => rxCsumVld,
        CSUM      => rxCsum
        );
  end generate INCLUDE_RX_CSUM;

  EXCLUDE_RX_CSUM: if (not (C_RXCSUM = 1)) generate
  begin
    rxCsum <= (others => '0');
    rxCsumVld <= '0';
  end generate EXCLUDE_RX_CSUM;

  -------------------------------------------------------------------------
  -- save partial csum value once calculated
  -------------------------------------------------------------------------

  SAVE_PARTIAL_CSUM_VAL : process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        raw_checksum <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (eof_reset = '1') then -- clear at end of frame
            raw_checksum <= (others => '0');
          elsif (rxCsumVld = '1') then
            raw_checksum <= rxCsum;
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- capture the statistics which is different for soft and hard TEMAC
  -------------------------------------------------------------------------

    frame_drop <= (EMAC_CLIENT_RX_STATS_VLD and not (rx_statistics_vector(27)));

    CAPTURE_STATS : process (RX_CLIENT_CLK)
    begin
      if rising_edge(RX_CLIENT_CLK) then
        if RESET2RX_CLIENT = '1' then
          statistics_vector <= (others => '0');
        else
          if (RX_CLIENT_CLK_ENBL = '1') then
            if (EMAC_CLIENT_RX_STATS_VLD = '1') then
              statistics_vector(25 downto 22) <= rx_statistics_vector(26 downto 23);
              statistics_vector(21 downto 0) <= rx_statistics_vector(21 downto 0);
            end if;
          end if;
        end if;
      end if;
    end process;



  -------------------------------------------------------------------------
  -- count the number of bytes in the frame being received for 8 bit interface
  -------------------------------------------------------------------------

  COUNT_FRAME_RX_BYTES : process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        frame_length_bytes <= (others => '0');
        frame_length_bytes_lat <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (end_of_frame_array(2) = '1') then -- clear at end of frame
            frame_length_bytes <= (others => '0');
          elsif (EMAC_CLIENT_RXD_VLD_LEGACY = '1') then
            frame_length_bytes <= frame_length_bytes + 1;
          end if;
          if (end_of_frame_array(2) = '1') then
            frame_length_bytes_lat <= frame_length_bytes;
          end if;	  
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- save the indication that we had a word 4 vlan tag strip
  -------------------------------------------------------------------------

  SAVE_WORD4_STRIP : process(RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        saveStripWord4VlanTag   <= '0';
      else
        if (stripWord4VlanTag = '1') then
              saveStripWord4VlanTag <= '1';
        elsif (end_of_frame_reset_in = '1') then
          saveStripWord4VlanTag <= '0';
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- save the indication that we had a word 4 vlan tag insertion
  -------------------------------------------------------------------------

  SAVE_WORD4_INSERT : process(RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        saveAutoInsertWord4VlanTag   <= '0';
      else
        if (autoInsertWord4VlanTag = '1') then
              saveAutoInsertWord4VlanTag <= '1';
        elsif (end_of_frame_reset_in = '1') then
          saveAutoInsertWord4VlanTag <= '0';
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- save the indication that we had a word 5 vlan tag insertion
  -------------------------------------------------------------------------

  SAVE_WORD5_INSERT : process(RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        saveAutoInsertWord5VlanTag   <= '0';
      else
        if (autoInsertWord5VlanTag = '1') then
              saveAutoInsertWord5VlanTag <= '1';
        elsif (end_of_frame_reset_in = '1') then
          saveAutoInsertWord5VlanTag <= '0';
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- save the good frame pulse so we can check it later
  -------------------------------------------------------------------------

  SAVE_GOOD_FRAME : process(RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        save_rx_goodframe   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (EMAC_CLIENT_RX_GOODFRAME_LEGACY = '1') then
                save_rx_goodframe <= '1';
          elsif (eof_reset = '1') then
            save_rx_goodframe <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- save the bad frame pulse so we can check it later
  -------------------------------------------------------------------------

  SAVE_BAD_FRAME : process(RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        save_rx_badframe   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (EMAC_CLIENT_RX_BADFRAME_LEGACY = '1') then
                save_rx_badframe <= '1';
          elsif (eof_reset = '1') then
            save_rx_badframe <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- check for not enough rxs memory
  -------------------------------------------------------------------------

  CHECK_RXS_MEM_AVAIL : process(RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        not_enough_rxs_memory   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          -- rxs_mem_last_read_out_ptr_cmb being read out of rxs memory during state END_OF_FRAME_CHECK_GOOD_BAD
          if (rxs_mem_addr_cntr   = unsigned(rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0)) or
              rxs_mem_addr_cntr+1 = unsigned(rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0)) or
              rxs_mem_addr_cntr+2 = unsigned(rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0)) or
              rxs_mem_addr_cntr+3 = unsigned(rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0)) or
              rxs_mem_addr_cntr+4 = unsigned(rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0)) or
              rxs_mem_addr_cntr+5 = unsigned(rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0))) then
                not_enough_rxs_memory <= '1';
          else
            not_enough_rxs_memory <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- create a pipeline of receive data, receive data valid, start of frame
  -- end of frame
  -------------------------------------------------------------------------

  PIPE_RX_INPUTS : process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        rx_data_words_array   <= (others => (others => '0'));
        rx_data_valid_array   <= (others => (others => '0'));
        rx_data_packed_ready_array <= (others => '0');
        start_of_frame_d1     <= '0';
        start_of_frame_array  <= (others => '0');
        end_of_frame_array    <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          rx_data_packed_ready_array (1) <= rx_data_packed_ready;
          if (rx_data_packed_ready = '1') then
            rx_data_words_array (1)     <= rx_data_packed_word;
            rx_data_valid_array (1)     <= rx_data_vld_packed_word;
          end if;
          start_of_frame_d1           <= EMAC_CLIENT_RXD_VLD_LEGACY;
          start_of_frame_array (1)    <= EMAC_CLIENT_RXD_VLD_LEGACY and not(start_of_frame_d1);
          end_of_frame_array (1)      <= start_of_frame_d1 and not(EMAC_CLIENT_RXD_VLD_LEGACY);
          for i in 1 to 7 loop
            rx_data_packed_ready_array (i+1)  <= rx_data_packed_ready_array (i);
            if (rx_data_packed_ready_array (i) = '1') then
              rx_data_words_array (i+1)  <= rx_data_words_array (i);
              rx_data_valid_array (i+1)  <= rx_data_valid_array (i);
            end if;
          end loop;
          for i in 1 to 28 loop
            start_of_frame_array (i+1)   <= start_of_frame_array (i);
          end loop;
          for i in 1 to 4 loop
            end_of_frame_array (i+1)     <= end_of_frame_array (i);
          end loop;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the destination address is broadcast
  -------------------------------------------------------------------------

  DETECT_BROADCAST : process(RX_CLIENT_CLK) -- valid by byte 10
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        frame_is_broadcast_d10   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (rx_data_words_array(1)(15 downto 0)  = X"FFFF" and
              rx_data_words_array(2)(31 downto 0) = X"FFFFFFFF" and
              start_of_frame_array(9) = '1') then
                frame_is_broadcast_d10 <= '1';
          elsif (eof_reset = '1') then
            frame_is_broadcast_d10 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the destination address is IP multicast
  -------------------------------------------------------------------------

  DETECT_IP_MULTICAST : process(RX_CLIENT_CLK) -- valid by byte 4
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        frame_is_ip_multicast_d4   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (rx_data_packed_word(31 downto 24) = X"5E" and
              rx_data_packed_word(23 downto 16) = X"00" and
              rx_data_packed_word(15 downto 8)  = X"01" and
              start_of_frame_array(3) = '1') then
                frame_is_ip_multicast_d4 <= '1';
          elsif (eof_reset = '1') then
            frame_is_ip_multicast_d4 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the destination address is any multicast
  -------------------------------------------------------------------------

  DETECT_MULTICAST : process(RX_CLIENT_CLK) -- valid by byte 10
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        frame_is_multicast_d10   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (rx_data_words_array(2)(0) = '1' and
              not((rx_data_words_array(1)(15 downto 0)  = X"FFFF")and
                  (rx_data_words_array(2)(31 downto 0) = X"FFFFFFFF"))and
              start_of_frame_array(9) = '1') then
                frame_is_multicast_d10 <= '1';
          elsif (eof_reset = '1') then
            frame_is_multicast_d10 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- save the destination (multicast) address for AXIStream status words
  -------------------------------------------------------------------------

  SAVE_DEST_ADDR : process(RX_CLIENT_CLK) -- valid by byte 10
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        multicast_addr_upper_d10   <= (others => '0');
        multicast_addr_lower_d10   <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (start_of_frame_array(9) = '1') then
            multicast_addr_upper_d10 <= rx_data_words_array(1)(15 downto 0);
            multicast_addr_lower_d10 <= rx_data_words_array(2)(31 downto 0);
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- save the bytes 12 thru 15 for AXIStream status words
  -------------------------------------------------------------------------

  SAVE_BYTES_12_TO_14 : process(RX_CLIENT_CLK) -- valid by byte 19
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        bytes_12_and_13_d19   <= (others => '0');
        bytes_14_and_15_d19   <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (start_of_frame_array(18) = '1') then
            bytes_12_and_13_d19 <= rx_data_words_array(1)(15 downto 0);
            bytes_14_and_15_d19 <= rx_data_words_array(1)(31 downto 16);
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame is a VLAN with type 8100
  -------------------------------------------------------------------------

  DETECT_VLAN_8100 : process(RX_CLIENT_CLK) -- valid by byte 15
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        frame_is_vlan_8100_d15   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = X"8100") and
              start_of_frame_array(14) = '1') then
                frame_is_vlan_8100_d15 <= '1';
          elsif (eof_reset = '1') then
            frame_is_vlan_8100_d15 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- Save the TPID value from the first VLAN tag
  -------------------------------------------------------------------------

  SAVE_FIRST_VLAN_TAG_VID : process(RX_CLIENT_CLK) -- valid by byte 17
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        first_vlan_tag_vid_d17   <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (start_of_frame_array(16) = '1') then
            first_vlan_tag_vid_d17 <= (rx_data_packed_word(19 downto 16) & rx_data_packed_word(31 downto 24));
          elsif (end_of_frame_reset_in = '1') then
            first_vlan_tag_vid_d17 <= (others => '0');
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- Save the TPID value from the second VLAN tag
  -------------------------------------------------------------------------

  SAVE_SECOND_VLAN_TAG_VID : process(RX_CLIENT_CLK) -- valid by byte 21
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        second_vlan_tag_vid_d21   <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (start_of_frame_array(20) = '1') then
            second_vlan_tag_vid_d21 <= (rx_data_packed_word(19 downto 16) & rx_data_packed_word(31 downto 24));
          elsif (end_of_frame_reset_in = '1') then
            second_vlan_tag_vid_d21 <= (others => '0');
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- Save the RX VLAN BRAM entry for the first VLAN tag TPID
  -------------------------------------------------------------------------

  SAVE_FIRST_VLAN_TAG_VID_BRAM_VALUE : process(RX_CLIENT_CLK) -- valid by byte 18
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        first_vlan_tag_bram_value_d18   <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (start_of_frame_array(17) = '1') then
            first_vlan_tag_bram_value_d18 <= RX_CL_CLK_VLAN_RD_DATA;
          elsif (end_of_frame_reset_in = '1') then
            first_vlan_tag_bram_value_d18 <= (others => '0');
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- Save the RX VLAN BRAM entry for the second VLAN tag TPID
  -------------------------------------------------------------------------

  SAVE_SECOND_VLAN_TAG_VID_BRAM_VALUE : process(RX_CLIENT_CLK) -- valid by byte 22
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        second_vlan_tag_bram_value_d22   <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (start_of_frame_array(21) = '1') then
            second_vlan_tag_bram_value_d22 <= RX_CL_CLK_VLAN_RD_DATA;
          elsif (end_of_frame_reset_in = '1') then
            second_vlan_tag_bram_value_d22 <= (others => '0');
          end if;
        end if;
      end if;
    end if;
  end process;

  RX_CL_CLK_VLAN_ADDR         <= (rx_data_packed_word(19 downto 16) & rx_data_packed_word(31 downto 24)) when (((start_of_frame_array(16) = '1') or (start_of_frame_array(20) = '1'))) else -- when RX_CL_CLK_VLAN_BRAM_EN_A = '1'
                                 rx_cl_clk_vlan_addr_reg; -- address stays the same to hold the value on the read output
  RX_CL_CLK_VLAN_BRAM_EN_A    <= '1' when ((start_of_frame_array(16) = '1') or (start_of_frame_array(20) = '1')) else
                                 '0';

  -------------------------------------------------------------------------
  -- don't allow the rx vlan addr to change when not reading to stabilize output
  -------------------------------------------------------------------------

  HOLD_RX_VLAN_ADDR : process(RX_CLIENT_CLK) -- valid by byte 15
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        rx_cl_clk_vlan_addr_reg   <= (others => '0');
      else
--        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((start_of_frame_array(16) = '1') or (start_of_frame_array(20) = '1'))) then                -- when RX_CL_CLK_VLAN_BRAM_EN_A = '1'
            rx_cl_clk_vlan_addr_reg <= (rx_data_packed_word(19 downto 16) & rx_data_packed_word(31 downto 24)); -- RX_CL_CLK_VLAN_ADDR store new address otherwise hold last address so read output stays the same while it is valid
          end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a first VLAN tag with type TPID 0
  -------------------------------------------------------------------------

  DETECT_FIRST_VLAN_TAG_TPID_0 : process(RX_CLIENT_CLK) -- valid by byte 15
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        first_tag_is_vlan_TPID_0_d15   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID0_REG_DATA(16 to 31)) and
              start_of_frame_array(14) = '1') then
                first_tag_is_vlan_TPID_0_d15 <= '1';
          elsif (eof_reset = '1') then
            first_tag_is_vlan_TPID_0_d15 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a first VLAN tag with type TPID 1
  -------------------------------------------------------------------------

  DETECT_FIRST_VLAN_TAG_TPID_1 : process(RX_CLIENT_CLK) -- valid by byte 15
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        first_tag_is_vlan_TPID_1_d15   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID0_REG_DATA(0 to 15)) and
              start_of_frame_array(14) = '1') then
                first_tag_is_vlan_TPID_1_d15 <= '1';
          elsif (eof_reset = '1') then
            first_tag_is_vlan_TPID_1_d15 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a first VLAN tag with type TPID 2
  -------------------------------------------------------------------------

  DETECT_FIRST_VLAN_TAG_TPID_2 : process(RX_CLIENT_CLK) -- valid by byte 15
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        first_tag_is_vlan_TPID_2_d15   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID1_REG_DATA(16 to 31)) and
              start_of_frame_array(14) = '1') then
                first_tag_is_vlan_TPID_2_d15 <= '1';
          elsif (eof_reset = '1') then
            first_tag_is_vlan_TPID_2_d15 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a first VLAN tag with type TPID 3
  -------------------------------------------------------------------------

  DETECT_FIRST_VLAN_TAG_TPID_3 : process(RX_CLIENT_CLK) -- valid by byte 15
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        first_tag_is_vlan_TPID_3_d15   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID1_REG_DATA(0 to 15)) and
              start_of_frame_array(14) = '1') then
                first_tag_is_vlan_TPID_3_d15 <= '1';
          elsif (eof_reset = '1') then
            first_tag_is_vlan_TPID_3_d15 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a second VLAN tag with type TPID 0
  -------------------------------------------------------------------------

  DETECT_SECOND_VLAN_TAG_TPID_0 : process(RX_CLIENT_CLK) -- valid by byte 19
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        second_tag_is_vlan_TPID_0_d19   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID0_REG_DATA(16 to 31)) and
              start_of_frame_array(18) = '1') then
                second_tag_is_vlan_TPID_0_d19 <= '1';
          elsif (eof_reset = '1') then
            second_tag_is_vlan_TPID_0_d19 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a second VLAN tag with type TPID 1
  -------------------------------------------------------------------------

  DETECT_SECOND_VLAN_TAG_TPID_1 : process(RX_CLIENT_CLK) -- valid by byte 19
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        second_tag_is_vlan_TPID_1_d19   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID0_REG_DATA(0 to 15)) and
              start_of_frame_array(18) = '1') then
                second_tag_is_vlan_TPID_1_d19 <= '1';
          elsif (eof_reset = '1') then
            second_tag_is_vlan_TPID_1_d19 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a second VLAN tag with type TPID 2
  -------------------------------------------------------------------------

  DETECT_SECOND_VLAN_TAG_TPID_2 : process(RX_CLIENT_CLK) -- valid by byte 19
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        second_tag_is_vlan_TPID_2_d19   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID1_REG_DATA(16 to 31)) and
              start_of_frame_array(18) = '1') then
                second_tag_is_vlan_TPID_2_d19 <= '1';
          elsif (eof_reset = '1') then
            second_tag_is_vlan_TPID_2_d19 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a second VLAN tag with type TPID 3
  -------------------------------------------------------------------------

  DETECT_SECOND_VLAN_TAG_TPID_3 : process(RX_CLIENT_CLK) -- valid by byte 19
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        second_tag_is_vlan_TPID_3_d19   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID1_REG_DATA(0 to 15)) and
              start_of_frame_array(18) = '1') then
                second_tag_is_vlan_TPID_3_d19 <= '1';
          elsif (eof_reset = '1') then
            second_tag_is_vlan_TPID_3_d19 <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame is a IPv4 Ethernet II frame with type 0800
  -------------------------------------------------------------------------

  DETECT_TYPE_0800 : process(RX_CLIENT_CLK) -- delay this check by one pipeline stage so we can detect vlan first valid by byte 22 when vlan
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        frame_has_type_0800_d22   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (frame_is_vlan_8100_d15 = '0') then -- no vlan
            if (((rx_data_words_array(1)(7 downto 0) & rx_data_words_array(1)(15 downto 8)) = X"0800") and start_of_frame_array(17) = '1') then
                    frame_has_type_0800_d22 <= '1';
            elsif (end_of_frame_reset_in = '1') then
              frame_has_type_0800_d22 <= '0';
            end if;
          else -- vlan
            if (((rx_data_words_array(1)(7 downto 0) & rx_data_words_array(1)(15 downto 8)) = X"0800") and start_of_frame_array(21) = '1') then
              frame_has_type_0800_d22 <= '1';
            elsif (end_of_frame_reset_in = '1') then
              frame_has_type_0800_d22 <= '0';
            end if;
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a valid length field
  -------------------------------------------------------------------------

  DETECT_VALID_LENGTH_FIELD : process(RX_CLIENT_CLK)-- delay this check by one pipeline stage so we can detect vlan first valid by byte 22 when vlan
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        frame_has_valid_length_field_d22   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (frame_is_vlan_8100_d15 = '0') then -- no vlan
            if (((rx_data_words_array(1)(7 downto 0) & rx_data_words_array(1)(15 downto 8)) < X"0601") and start_of_frame_array(17) = '1') then
              frame_has_valid_length_field_d22 <= '1';
            elsif (end_of_frame_reset_in = '1') then
              frame_has_valid_length_field_d22 <= '0';
            end if;
          else -- vlan
            if (((rx_data_words_array(1)(7 downto 0) & rx_data_words_array(1)(15 downto 8)) < X"0601") and start_of_frame_array(21) = '1') then
              frame_has_valid_length_field_d22 <= '1';
            elsif (end_of_frame_reset_in = '1') then
              frame_has_valid_length_field_d22 <= '0';
            end if;
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- detect if the frame is a IPv4 Ethernet SNAP frame with type 0800
  -------------------------------------------------------------------------

  DETECT_SNAP : process(RX_CLIENT_CLK)-- delay this check by one pipeline stage so we can detect vlan first valid by byte 30 when vlan
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        frame_is_snap_d30   <= '0';
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (frame_is_vlan_8100_d15 = '0') then -- no vlan
            if ((rx_data_words_array(3)(31 downto 16) = X"AAAA") and
                 (rx_data_words_array(2)(31 downto 0) =  X"00000003") and
                 (rx_data_words_array(1)(15 downto 0) =  X"0008") and
                 start_of_frame_array(25) = '1') and (frame_has_valid_length_field_d22 = '1') then
                   frame_is_snap_d30 <= '1';
            elsif (end_of_frame_reset_in = '1') then
              frame_is_snap_d30 <= '0';
            end if;
          else -- vlan
            if ((rx_data_words_array(3)(31 downto 16) = X"AAAA") and
                 (rx_data_words_array(2)(31 downto 0) =  X"00000003") and
                 (rx_data_words_array(1)(15 downto 0) =  X"0008") and
                 start_of_frame_array(29) = '1') and (frame_has_valid_length_field_d22 = '1') then
                   frame_is_snap_d30 <= '1';
            elsif (end_of_frame_reset_in = '1') then
              frame_is_snap_d30 <= '0';
            end if;
          end if;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- Initialize the dual port address for the RXD memory
  -------------------------------------------------------------------------
  RXD_ADDR_CNTR: process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        rxd_mem_addr_cntr  <= rxd_mem_empty_mask;
      elsif (rxd_addr_cntr_load = '1') then
        rxd_mem_addr_cntr  <= unsigned(rxd_mem_next_available4write_ptr_cmb);
      else
        if (rxd_addr_cntr_en = '1' and rx_data_packed_ready_array(3) = '1' and RX_CLIENT_CLK_ENBL = '1' and not(stripWord4VlanTag = '1')) then
          rxd_mem_addr_cntr  <= rxd_mem_addr_cntr + 1;
        elsif ((autoInsertWord4VlanTag = '1' or autoInsertWord5VlanTag = '1')and RX_CLIENT_CLK_ENBL = '1') then -- I think we need to check for RX_CLIENT_CLK_ENBL = '1' here
            rxd_mem_addr_cntr  <= rxd_mem_addr_cntr + 1;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- Initialize the dual port address for the RXS memory
  -------------------------------------------------------------------------
  RXS_ADDR_CNTR: process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        rxs_mem_addr_cntr  <= rxs_mem_four_mask;
      elsif (rxs_addr_cntr_load = '1') then
        rxs_mem_addr_cntr  <= unsigned(rxs_mem_next_available4write_ptr_cmb);
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          if (rxs_addr_cntr_en = '1' and not(rxs_mem_addr_cntr = rxs_mem_full_mask)) then
            rxs_mem_addr_cntr  <= rxs_mem_addr_cntr + 1;
          elsif (rxs_addr_cntr_en = '1' and rxs_mem_addr_cntr = rxs_mem_full_mask) then
            rxs_mem_addr_cntr  <= rxs_mem_four_mask;
          end if;
        end if;
      end if;
    end if;
  end process;

  RX_CLIENT_RXS_DPMEM_ADDR(C_RXS_MEM_ADDR_WIDTH downto 0) <=
    std_logic_vector(rxs_mem_one_mask)   when receive_frame_current_state = RESET_INIT_MEM_PTR_2 else
    std_logic_vector(rxs_mem_two_mask)   when receive_frame_current_state = RESET_INIT_MEM_PTR_3 else
    std_logic_vector(rxs_mem_three_mask) when receive_frame_current_state = RESET_INIT_MEM_PTR_4 else
    std_logic_vector(rxs_mem_two_mask)   when receive_frame_current_state = UPDATE_MEM_PTR_2 else
    std_logic_vector(rxs_mem_addr_cntr);

  RX_CLIENT_RXS_DPMEM_WR_EN(0) <=
    '1'  when receive_frame_current_state = RESET_INIT_MEM_PTR_2 else
    '1'  when receive_frame_current_state = RESET_INIT_MEM_PTR_3 else
    '1'  when receive_frame_current_state = RESET_INIT_MEM_PTR_4 else
    '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_1 else
    '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_2 else
    '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_3 else
    '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_4 else
    '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_5 else
    '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_6 else
    '1'  when receive_frame_current_state = UPDATE_MEM_PTR_2 else
    '0';

  RX_CLIENT_RXS_DPMEM_WR_DATA(35 downto 0) <=
    zero_extend_rxd_mask36 & rxd_mem_last_read_out_ptr_cmb        when receive_frame_current_state = RESET_INIT_MEM_PTR_2 else
    zero_extend_rxs_mask36 & rxs_mem_next_available4write_ptr_cmb when receive_frame_current_state = RESET_INIT_MEM_PTR_3 else
    zero_extend_rxs_mask36 & std_logic_vector(rxs_mem_full_mask)  when receive_frame_current_state = RESET_INIT_MEM_PTR_4 else
    zero_extend_rxs_mask36 & rxs_mem_next_available4write_ptr_cmb when receive_frame_current_state = UPDATE_MEM_PTR_2 else
    rxs_status_word_1_cmb                                         when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_1 else
    rxs_status_word_2                                         when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_2 else
    rxs_status_word_3                                         when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_3 else
    rxs_status_word_4                                         when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_4 else
    rxs_status_word_5                                         when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_5 else
    rxs_status_word_6_cmb                                     when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_6 else
    (others => '0');

  RX_CLIENT_RXD_DPMEM_WR_EN(0) <=
    '1'                           when autoInsertWord4VlanTag = '1' else -- tag before word 4
    '1'                           when autoInsertWord5VlanTag = '1' else -- tag before word 5 (word 4 was stripped)
    rx_data_packed_ready_array(3) when receive_frame_data_current_state = RECEIVING_FRAME and not(stripWord4VlanTag = '1') else -- normal and block when stripping word 4
    '0';

  autoInsertWord4VlanTag <= '1' when word4TagEnabled_d18 = '1'   and start_of_frame_array(18) = '1' else -- tag before word 4
                            '0';
  autoInsertWord5VlanTag <= '1' when word5TagEnabled_d22 = '1'   and start_of_frame_array(22) = '1' else -- tag before word 5 (word 4 was stripped)
                            '0';
  translateWord4VlanVid  <= '1' when word4TransEnabled_d18 = '1' and start_of_frame_array(19) = '1' else -- translate word 4 VID
                            '0';
  translateWord5VlanVid  <= '1' when word5TransEnabled_d19 = '1' and start_of_frame_array(23) = '1' else -- translate word 5 VID
                            '0';
  stripWord4VlanTag      <= '1' when word4StrpEnabled_d18 = '1'  and start_of_frame_array(19) = '1' else -- stripping word 4
                            '0';
  --------------------------------------------------------------------------
  -- when stripping and tagging we need to adjust byte count and adjust RXD
  -- address counter
  --------------------------------------------------------------------------

  RX_CLIENT_RXD_DPMEM_ADDR(C_RXD_MEM_ADDR_WIDTH downto 0) <= std_logic_vector(rxd_mem_addr_cntr);

  RX_CLIENT_RXD_DPMEM_WR_DATA(35 downto 0) <=
    X"f" & RX_CL_CLK_RX_TAG_REG_DATA(24 to 31) & RX_CL_CLK_RX_TAG_REG_DATA(16 to 23) & RX_CL_CLK_RX_TAG_REG_DATA(8 to 15) & RX_CL_CLK_RX_TAG_REG_DATA(0 to 7) when autoInsertWord4VlanTag = '1' else -- tag before word 4
    X"f" & RX_CL_CLK_RX_TAG_REG_DATA(24 to 31) & RX_CL_CLK_RX_TAG_REG_DATA(16 to 23) & RX_CL_CLK_RX_TAG_REG_DATA(8 to 15) & RX_CL_CLK_RX_TAG_REG_DATA(0 to 7) when autoInsertWord5VlanTag = '1' else -- tag before word 5 (word 4 was stripped)
    X"f" & first_vlan_tag_bram_value_d18(22 to 29)  & rx_data_words_array(2)(23 downto 20) & first_vlan_tag_bram_value_d18(18 to 21)  & rx_data_words_array(2)(15 downto 0) when  translateWord4VlanVid = '1' else -- translate word 4 VID
    X"f" & second_vlan_tag_bram_value_d22(22 to 29) & rx_data_words_array(2)(23 downto 20) & second_vlan_tag_bram_value_d22(18 to 21) & rx_data_words_array(2)(15 downto 0) when  translateWord5VlanVid = '1' else -- translate word 5 VID
    rx_data_valid_array(2) & rx_data_words_array(2); -- normal case

  --------------------------------------------------------------------------
  -- receive frame State Machine
  -- RXFRMSM_REGS_PROCESS: registered process of the state machine
  -- RXFRMSM_CMB_PROCESS:  combinatorial next-state logic
  --------------------------------------------------------------------------

  RXFRMSM_REGS_PROCESS: process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        receive_frame_current_state          <= RESET_INIT_MEM_PTR_1;
        receive_frame_data_current_state     <= RESET;	
        rxd_mem_next_available4write_ptr_reg <= std_logic_vector(rxd_mem_empty_mask);
        rxd_mem_last_read_out_ptr_reg        <= std_logic_vector(rxd_mem_full_mask);
        rxs_mem_next_available4write_ptr_reg <= std_logic_vector(rxs_mem_four_mask);
        rxs_status_word_1_reg                <= (others => '0');
        rxs_status_word_6_reg                <= (others => '0');
      else
        if (RX_CLIENT_CLK_ENBL = '1') then
          receive_frame_current_state          <= receive_frame_next_state;
          receive_frame_data_current_state     <= receive_frame_data_next_state;	  
          rxd_mem_next_available4write_ptr_reg <= rxd_mem_next_available4write_ptr_cmb;
          rxd_mem_last_read_out_ptr_reg        <= rxd_mem_last_read_out_ptr_cmb;
          rxs_mem_next_available4write_ptr_reg <= rxs_mem_next_available4write_ptr_cmb;
          rxs_status_word_1_reg                <= rxs_status_word_1_cmb;
          rxs_status_word_6_reg                <= rxs_status_word_6_cmb;
        end if;
      end if;
    end if;
  end process;


  RX_RECEIVEFSM_CMD_PROCESS: process (
    receive_frame_data_current_state,
    start_of_frame_array,
    end_of_frame_array,
    save_rx_goodframe,
    save_rx_badframe,
    rxd_mem_next_available4write_ptr_reg,
    rxd_mem_next_available4write_ptr_cmb,
    rx_data_packed_ready,
    rxd_mem_last_read_out_ptr_reg,
    rxd_mem_last_read_out_ptr_cmb,
    rxs_status_word_1_reg,
    rxs_status_word_1_cmb,
    rxs_status_word_6_reg,
    rxs_status_word_6_cmb,
    rxd_mem_addr_cntr,
    not_enough_rxs_memory,
    RX_CL_CLK_BRDCAST_REJ,
    RX_CL_CLK_MULCAST_REJ,
    frame_is_broadcast_d10,
    frame_is_multicast_d10,
    saveExtendedMulticastReject,
    rxd_mem_empty_mask,
    rxd_mem_full_mask,
    rxclclk_rxd_mem_last_read_out_ptr_d1,
    frame_length_bytes_lat,
    saveAutoInsertWord4VlanTag,
    saveStripWord4VlanTag,
    saveAutoInsertWord5VlanTag,
    RX_CL_CLK_BAD_FRAME_ENBL
    )
  begin

    rxd_addr_cntr_en              <= '0';
    rxd_addr_cntr_load            <= '0';
    RX_FRAME_RECEIVED_INTRPT      <= '0';
    RX_FRAME_REJECTED_INTRPT      <= '0';
    RX_BUFFER_MEM_OVERFLOW_INTRPT <= '0';
    update_status_fifo            <= '0';

    rxd_mem_next_available4write_ptr_cmb <= rxd_mem_next_available4write_ptr_reg;
    rxd_mem_last_read_out_ptr_cmb        <= rxd_mem_last_read_out_ptr_reg;
    rxs_status_word_1_cmb                <= rxs_status_word_1_reg;
    rxs_status_word_6_cmb(15 downto 0)   <= rxs_status_word_6_reg(15 downto 0);

    case receive_frame_data_current_state is

      when RESET =>
              receive_frame_data_next_state        <= WAIT_FOR_START_OF_FRAME;
        rxd_mem_next_available4write_ptr_cmb <= std_logic_vector(rxd_mem_empty_mask);
        rxd_mem_last_read_out_ptr_cmb        <= std_logic_vector(rxd_mem_full_mask);
        rxs_status_word_1_cmb                <= (others => '0');

      when WAIT_FOR_START_OF_FRAME =>
        rxd_mem_last_read_out_ptr_cmb    <= rxclclk_rxd_mem_last_read_out_ptr_d1(C_RXD_MEM_ADDR_WIDTH downto 0);
        rxd_addr_cntr_load               <= '1';
        if (start_of_frame_array (5) = '1') then
          receive_frame_data_next_state  <= RECEIVING_FRAME;
        else
          receive_frame_data_next_state  <= WAIT_FOR_START_OF_FRAME;
        end if;

      when RECEIVING_FRAME =>
        rxd_mem_last_read_out_ptr_cmb    <= rxclclk_rxd_mem_last_read_out_ptr_d1(C_RXD_MEM_ADDR_WIDTH downto 0);
        rxs_status_word_1_cmb(15 downto C_RXD_MEM_ADDR_WIDTH+1) <= (others => '0');
        rxs_status_word_1_cmb(C_RXD_MEM_ADDR_WIDTH downto 0)    <= rxd_mem_next_available4write_ptr_cmb;
        rxd_addr_cntr_en                 <= '1';
        if (std_logic_vector(rxd_mem_addr_cntr) = rxd_mem_last_read_out_ptr_cmb and rx_data_packed_ready = '1') then -- RXD memory overflow
          receive_frame_data_next_state  <= WAIT_FOR_START_OF_FRAME;
          RX_BUFFER_MEM_OVERFLOW_INTRPT  <= '1';
        elsif (end_of_frame_array (5) = '0') then
          receive_frame_data_next_state  <= RECEIVING_FRAME;
        else
          receive_frame_data_next_state  <= END_OF_FRAME_CHECK_GOOD_BAD;
        end if;

      when END_OF_FRAME_CHECK_GOOD_BAD =>
        rxs_status_word_1_cmb(35 downto 32)  <= (others => '0');
        if (saveAutoInsertWord4VlanTag = '1' and saveStripWord4VlanTag = '0') then
          rxs_status_word_1_cmb(31 downto 16)  <= std_logic_vector(frame_length_bytes_lat + 4);
          rxs_status_word_6_cmb(15 downto 0)   <= std_logic_vector(frame_length_bytes_lat + 4);
        elsif (saveStripWord4VlanTag = '1' and saveAutoInsertWord5VlanTag = '0' and saveAutoInsertWord4VlanTag = '0') then
          rxs_status_word_1_cmb(31 downto 16)  <= std_logic_vector(frame_length_bytes_lat - 4);
          rxs_status_word_6_cmb(15 downto 0)   <= std_logic_vector(frame_length_bytes_lat - 4);
        else
          rxs_status_word_1_cmb(31 downto 16)  <= std_logic_vector(frame_length_bytes_lat);
          rxs_status_word_6_cmb(15 downto 0)   <= std_logic_vector(frame_length_bytes_lat);
        end if;
        if (not_enough_rxs_memory = '1') then  -- RXS memory overflow
          receive_frame_data_next_state       <= WAIT_FOR_START_OF_FRAME;
          RX_BUFFER_MEM_OVERFLOW_INTRPT  <= '1';
        elsif ((save_rx_goodframe = '1') or (save_rx_badframe = '1' and RX_CL_CLK_BAD_FRAME_ENBL = '1'))  then
          if ((frame_is_broadcast_d10 = '1' and RX_CL_CLK_BRDCAST_REJ = '1') or
              (frame_is_multicast_d10 = '1' and RX_CL_CLK_MULCAST_REJ = '1') or
              (saveExtendedMulticastReject = '1'))then
            receive_frame_data_next_state       <= WAIT_FOR_START_OF_FRAME;
            RX_FRAME_REJECTED_INTRPT     <= '1';
          else
            rxd_mem_next_available4write_ptr_cmb <= std_logic_vector(rxd_mem_addr_cntr);
            update_status_fifo           <= '1';	    
            receive_frame_data_next_state       <= WAIT_FOR_START_OF_FRAME;
            RX_FRAME_RECEIVED_INTRPT     <= '1';
          end if;
        elsif (save_rx_badframe = '1') then
          receive_frame_data_next_state       <= WAIT_FOR_START_OF_FRAME;
          RX_FRAME_REJECTED_INTRPT       <= '1';
        else
          receive_frame_data_next_state  <= END_OF_FRAME_CHECK_GOOD_BAD;
        end if;

      when others   =>
        receive_frame_data_next_state    <= WAIT_FOR_START_OF_FRAME;
    end case;
  end process;



  RXFRMSM_CMB_PROCESS : process (
    receive_frame_current_state,
    rxs_mem_addr_cntr,
    rxs_mem_next_available4write_ptr_cmb,
    update_status_fifo, rxs_mem_next_available4write_ptr_reg,
    rxs_mem_four_mask
    )
  begin

    rxs_addr_cntr_en              <= '0';
    rxs_addr_cntr_load            <= '0';
    rxs_mem_next_available4write_ptr_cmb <= rxs_mem_next_available4write_ptr_reg;

    case receive_frame_current_state is

      when RESET_INIT_MEM_PTR_1 =>
        receive_frame_next_state             <= RESET_INIT_MEM_PTR_2;
        rxs_mem_next_available4write_ptr_cmb <= std_logic_vector(rxs_mem_four_mask);

      when RESET_INIT_MEM_PTR_2 =>
        receive_frame_next_state         <= RESET_INIT_MEM_PTR_3;

      when RESET_INIT_MEM_PTR_3 =>
        receive_frame_next_state         <= RESET_INIT_MEM_PTR_4;

      when RESET_INIT_MEM_PTR_4 =>
        receive_frame_next_state         <= IDLE;

      when IDLE => 
          if (update_status_fifo = '1') then
              receive_frame_next_state   <= UPDATE_STATUS_FIFO_WORD_1;
          else
              receive_frame_next_state   <= IDLE;
          end if;
          rxs_addr_cntr_load             <= '1';

      when UPDATE_STATUS_FIFO_WORD_1 =>
        receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_2;
        rxs_addr_cntr_en                 <= '1';

      when UPDATE_STATUS_FIFO_WORD_2 =>
        receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_3;
        rxs_addr_cntr_en                 <= '1';

      when UPDATE_STATUS_FIFO_WORD_3 =>
        receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_4;
        rxs_addr_cntr_en                 <= '1';

      when UPDATE_STATUS_FIFO_WORD_4 =>
        receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_5;
        rxs_addr_cntr_en                 <= '1';

      when UPDATE_STATUS_FIFO_WORD_5 =>
        receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_6;
        rxs_addr_cntr_en                 <= '1';

      when UPDATE_STATUS_FIFO_WORD_6 =>
        receive_frame_next_state         <= UPDATE_MEM_PTR_1;
        rxs_addr_cntr_en                 <= '1';

      when UPDATE_MEM_PTR_1 =>
        receive_frame_next_state         <= UPDATE_MEM_PTR_2;
        rxs_mem_next_available4write_ptr_cmb <= std_logic_vector(rxs_mem_addr_cntr);

      when UPDATE_MEM_PTR_2 =>
              receive_frame_next_state         <= IDLE;

      when others   =>
        receive_frame_next_state         <= RESET_INIT_MEM_PTR_1;
    end case;
  end process;

  -------------------------------------------------------------------------
  -- check enhanced multicast address filtering or not
  -------------------------------------------------------------------------

  EXTENDED_MULTICAST: if(C_MCAST_EXTEND = 1) generate

    type EMCFLTRSM_TYPE is (
      WAIT_FRAME_START,
      GET_SECOND_BYTE,
      GET_THIRD_BYTE,
      GET_FORTH_BYTE,
      GET_FIFTH_BYTE,
      READ_TABLE_ENTRY,
      READ_TABLE_ENTRY2,
      GET_UNI_ADDRESS,
      CHECK_UNI_ADDRESS,
      GET_BRDCAST_ADDRESS,
      CHECK_BRDCAST_ADDRESS,
      ACCEPT_AND_WAIT_TILL_END,
      REJECT_AND_WAIT_TILL_END
    );

    signal eMcFltrSM_Cs           : EMCFLTRSM_TYPE;
    signal eMcFltrSM_Ns           : EMCFLTRSM_TYPE;
    signal tempDestAddr           : std_logic_vector(0 to 47);
    signal unicastMatch           : std_logic;
    signal broadcastMatch         : std_logic;
    signal emacClientRxdLegacy_d1 : std_logic_vector(7 downto 0);

    signal rxClClkMcastEn_i        : std_logic;
    signal rxClClkMcastAddr_i      : std_logic_vector(0 to 14);
    signal rxClClkMcastAddr_i_d    : std_logic_vector(0 to 14);
    signal rx_cl_clk_mcast_rd_data_d1 : std_logic;

  begin

  RX_CL_CLK_MCAST_EN   <= rxClClkMcastEn_i;
  RX_CL_CLK_MCAST_ADDR <= rxClClkMcastAddr_i;

    process(RX_CLIENT_CLK)
      begin
        if(rising_edge(RX_CLIENT_CLK)) then
          if(RESET2RX_CLIENT='1') then
            emacClientRxdLegacy_d1     <= (others => '0');
            rx_cl_clk_mcast_rd_data_d1 <= '0';
          else
            rx_cl_clk_mcast_rd_data_d1 <= RX_CL_CLK_MCAST_RD_DATA(0);
            if(RX_CLIENT_CLK_ENBL='1') then
              emacClientRxdLegacy_d1   <= EMAC_CLIENT_RXD_LEGACY;
            end if;
          end if;
        end if;
    end process;

    COMPARE_UNICAST_ADDR_PROCESS: process (RX_CLIENT_CLK)
    begin
      if (RX_CLIENT_CLK'event and RX_CLIENT_CLK = '1') then
        if (RESET2RX_CLIENT = '1') then
          unicastMatch <= '0';
        else
          if (tempDestAddr(0 to 7)   = RX_CL_CLK_UAWL_REG_DATA(24 to 31) and
              tempDestAddr(8 to 15)  = RX_CL_CLK_UAWL_REG_DATA(16 to 23) and
              tempDestAddr(16 to 23) = RX_CL_CLK_UAWL_REG_DATA(8 to 15) and
              tempDestAddr(24 to 31) = RX_CL_CLK_UAWL_REG_DATA(0 to 7) and
              tempDestAddr(32 to 39) = RX_CL_CLK_UAWU_REG_DATA(24 to 31) and
              tempDestAddr(40 to 47) = RX_CL_CLK_UAWU_REG_DATA(16 to 23))then
            unicastMatch <= '1';
          else
            unicastMatch <= '0';
          end if;
        end if;
      end if;
    end process;

    COMPARE_BROADCAST_ADDR_PROCESS: process (RX_CLIENT_CLK)
    begin
      if (RX_CLIENT_CLK'event and RX_CLIENT_CLK = '1') then
        if (RESET2RX_CLIENT = '1') then
          broadcastMatch <= '0';
        else
          if (tempDestAddr=x"ffffffffffff") then
            broadcastMatch <= '1';
          else
            broadcastMatch <= '0';
          end if;
        end if;
      end if;
    end process;

    CAPTURE_TEMPDESTADDR_PROCESS: process (RX_CLIENT_CLK)
    begin
      if (RX_CLIENT_CLK'event and RX_CLIENT_CLK = '1') then
        if (RESET2RX_CLIENT = '1') then
          tempDestAddr    <= (others => '0');
        else
          if (RX_CLIENT_CLK_ENBL = '1') then
            if (start_of_frame_array (1) = '1') then
              tempDestAddr(0 to 7)   <= emacClientRxdLegacy_d1(7 downto 0);
              tempDestAddr(8 to 47)  <= (others => '0');
            elsif (start_of_frame_array (2) = '1') then
              tempDestAddr(0 to 7)   <= tempDestAddr(0 to 7);
              tempDestAddr(8 to 15)  <= emacClientRxdLegacy_d1(7 downto 0);
              tempDestAddr(16 to 47) <= (others => '0');
            elsif (start_of_frame_array (3) = '1') then
              tempDestAddr(0 to 15)  <= tempDestAddr(0 to 15);
              tempDestAddr(16 to 23) <= emacClientRxdLegacy_d1(7 downto 0);
              tempDestAddr(24 to 47) <= (others => '0');
            elsif (start_of_frame_array (4) = '1') then
              tempDestAddr(0 to 23)  <= tempDestAddr(0 to 23);
              tempDestAddr(24 to 31) <= emacClientRxdLegacy_d1(7 downto 0);
              tempDestAddr(32 to 47) <= (others => '0');
            elsif (start_of_frame_array (5) = '1') then
              tempDestAddr(0 to 31)  <= tempDestAddr(0 to 31);
              tempDestAddr(32 to 39) <= emacClientRxdLegacy_d1(7 downto 0);
              tempDestAddr(40 to 47) <= (others => '0');
            elsif (start_of_frame_array (6) = '1') then
              tempDestAddr(0 to 39)  <= tempDestAddr(0 to 39);
              tempDestAddr(40 to 47) <= emacClientRxdLegacy_d1(7 downto 0);
            else
              tempDestAddr(0 to 47)  <= tempDestAddr(0 to 47);
            end if;
          end if;
        end if;
      end if;
    end process;

  -------------------------------------------------------------------------
  -- save the indication that we had an extended multicast reject
  -------------------------------------------------------------------------

  SAVE_EXTENDED_MULTICAST_REJECT : process(RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        saveExtendedMulticastReject   <= '0';
      else
        if (eof_reset = '1') then
          saveExtendedMulticastReject <= '0';
        elsif (extendedMulticastReject = '1') then
              saveExtendedMulticastReject <= '1';
        end if;
      end if;
    end if;
  end process;

    EMCFLTRSM_REGS_PROCESS: process (RX_CLIENT_CLK )
    begin
      if (RX_CLIENT_CLK'event and RX_CLIENT_CLK = '1') then
        if (RESET2RX_CLIENT = '1') then
          eMcFltrSM_Cs     <= WAIT_FRAME_START;
          rxClClkMcastAddr_i_d <= (others => '0');
        else
          if (RX_CLIENT_CLK_ENBL = '1') then
            eMcFltrSM_Cs <= eMcFltrSM_Ns;
            rxClClkMcastAddr_i_d <= rxClClkMcastAddr_i;
          end if;
        end if;
      end if;
    end process;

    EMCFLTRSM_CMB_PROCESS: process (
       eMcFltrSM_Cs,
       start_of_frame_array (1),
       end_of_frame_array (1),
       RX_CL_CLK_NEW_FNC_ENBL,
       RX_CL_CLK_EMULTI_FLTR_ENBL,
       emacClientRxdLegacy_d1,
       RX_CL_CLK_MCAST_RD_DATA,
       rx_cl_clk_mcast_rd_data_d1,
       tempDestAddr,
       RX_CL_CLK_UAWL_REG_DATA,
       RX_CL_CLK_UAWU_REG_DATA,
       start_of_frame_array (8),
       unicastMatch,
       rxClClkMcastAddr_i_d,
       rxClClkMcastAddr_i,
       broadcastMatch,
       eof_reset
     )
    begin

      extendedMulticastReject   <= '0';
      rxClClkMcastEn_i          <= '0';
      rxClClkMcastAddr_i        <= rxClClkMcastAddr_i_d;

      case eMcFltrSM_Cs is

        when WAIT_FRAME_START =>
          rxClClkMcastAddr_i <= (others => '0');
          if (RX_CL_CLK_NEW_FNC_ENBL = '1' and RX_CL_CLK_EMULTI_FLTR_ENBL = '1') then
            if (start_of_frame_array (1) = '1')then
              if (emacClientRxdLegacy_d1=X"01")then
                eMcFltrSM_Ns <= GET_SECOND_BYTE; -- looks like IP generated multicast so far
              elsif (emacClientRxdLegacy_d1(0)='0')then
                eMcFltrSM_Ns <= GET_UNI_ADDRESS; -- it's a unicast address that we need to compare
              elsif (emacClientRxdLegacy_d1=X"FF")then
                eMcFltrSM_Ns <= GET_BRDCAST_ADDRESS; -- looks like broadcast so far
              else
                eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END; -- must be multicast but non-IP generated
                extendedMulticastReject <= '1';
              end if;
            else
              eMcFltrSM_Ns <= WAIT_FRAME_START; -- a new frame hasn't started yet
            end if;
          else
            eMcFltrSM_Ns <= WAIT_FRAME_START; -- extended multicast filtering not enabled
          end if;

        when GET_SECOND_BYTE =>
          if (emacClientRxdLegacy_d1=X"00")then
            eMcFltrSM_Ns <= GET_THIRD_BYTE; -- still looks like IP generated multicast so far
          else
            eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END; -- must be multicast but non-IP generated
            extendedMulticastReject <= '1';
          end if;

        when GET_THIRD_BYTE =>
          if (emacClientRxdLegacy_d1=X"5e")then
            eMcFltrSM_Ns <= GET_FORTH_BYTE; -- it is an IP generated multicast so let get the rest and look it up
          else
            eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END; -- must be multicast but non-IP generated
            extendedMulticastReject <= '1';
          end if;

        when GET_FORTH_BYTE =>
          rxClClkMcastAddr_i(0 to 6) <= emacClientRxdLegacy_d1(6 downto 0);
          eMcFltrSM_Ns <= GET_FIFTH_BYTE;

        when GET_FIFTH_BYTE =>
          rxClClkMcastAddr_i(7 to 14) <= emacClientRxdLegacy_d1(7 downto 0);
          rxClClkMcastEn_i            <= '1';
          eMcFltrSM_Ns <= READ_TABLE_ENTRY;

        when READ_TABLE_ENTRY =>
          --rxClClkMcastAddr_i(7 to 14) <= emacClientRxdLegacy_d1(7 downto 0);
          rxClClkMcastEn_i            <= '1';
          eMcFltrSM_Ns <= READ_TABLE_ENTRY2;

        when READ_TABLE_ENTRY2 =>
          rxClClkMcastEn_i            <= '1';
          if (rx_cl_clk_mcast_rd_data_d1 ='0')then
            eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END;
            extendedMulticastReject  <= '1';
          else
            eMcFltrSM_Ns <= ACCEPT_AND_WAIT_TILL_END;
          end if;

        when GET_UNI_ADDRESS =>
          if (start_of_frame_array (8)='1')then
            eMcFltrSM_Ns <= CHECK_UNI_ADDRESS;
          else
            eMcFltrSM_Ns <= GET_UNI_ADDRESS;
          end if;

        when GET_BRDCAST_ADDRESS =>
          if (start_of_frame_array (8)='1')then
            eMcFltrSM_Ns <= CHECK_BRDCAST_ADDRESS;
          else
            eMcFltrSM_Ns <= GET_BRDCAST_ADDRESS;
          end if;

        when CHECK_BRDCAST_ADDRESS =>
          if (broadcastMatch='1')then
            eMcFltrSM_Ns <= ACCEPT_AND_WAIT_TILL_END;
          else
            eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END;
            extendedMulticastReject  <= '1';
          end if;

        when CHECK_UNI_ADDRESS =>
          if (unicastMatch = '1')then
            eMcFltrSM_Ns <= ACCEPT_AND_WAIT_TILL_END;
          else
            eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END;
            extendedMulticastReject  <= '1';
          end if;

        when REJECT_AND_WAIT_TILL_END =>
          if (eof_reset = '1' )then
            eMcFltrSM_Ns <= WAIT_FRAME_START;
            extendedMulticastReject  <= '0';
          else
            eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END;
            extendedMulticastReject  <= '1';
          end if;

        when ACCEPT_AND_WAIT_TILL_END =>
          extendedMulticastReject  <= '0';
          if (eof_reset = '1' )then
            eMcFltrSM_Ns <= WAIT_FRAME_START;
          else
            eMcFltrSM_Ns <= ACCEPT_AND_WAIT_TILL_END;
          end if;

        when others   =>
          eMcFltrSM_Ns <= WAIT_FRAME_START;
      end case;
    end process;


  end generate EXTENDED_MULTICAST;

  NO_EXTENDED_MULTICAST: if(C_MCAST_EXTEND = 0) generate
  begin
    extendedMulticastReject <= '0';
    RX_CL_CLK_MCAST_ADDR    <= (others => '0');
    RX_CL_CLK_MCAST_EN      <= '0';
    saveExtendedMulticastReject <= '0';
  end generate NO_EXTENDED_MULTICAST;

end rtl;


------------------------------------------------------------------------------
-- rx_emac_if.vhd
------------------------------------------------------------------------------
-- (c) Copyright 2004-2009 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, rtlLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-- ------------------------------------------------------------------------------
--
------------------------------------------------------------------------------
-- Filename:        rx_emac_if.vhd
-- Version:         v1.00a
-- Description:     Receive interface between AXIStream and Temac
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to rtlrove
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:          MSH
--
--  MSH     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of : out   std_logic; port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Libraries used;
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.rx_if_pack.all;

library work;
use work.clock_cross_pack.all;

-------------------------------------------------------------------------------
-- Definition of Generics :
-------------------------------------------------------------------------------
-- System generics
--  C_FAMILY              -- Xilinx FPGA Family
--  C_RXD_MEM_BYTES               -- Depth of RX memory in Bytes
--  C_RXCSUM
--     0  No checksum offloading
--     1  Partial (legacy) checksum offloading
--     2  Full checksum offloading
--  C_RXVLAN_TRAN         -- Enable RX enhanced VLAN translation
--  C_RXVLAN_TAG          -- Enable RX enhanced VLAN taging
--  C_RXVLAN_STRP         -- Enable RX enhanced VLAN striping
--  C_MCAST_EXTEND        -- Enable RX extended multicast address filtering

-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Definition of Ports :
-------------------------------------------------------------------------------
--    BUS2IP_CLK
--    BUS2IP_RESET
--
--    AXI_STR_RXD_ACLK
--    AXI_STR_RXD_ARESET
--    AXI_STR_RXD_VALID
--    AXI_STR_RXD_READY
--    AXI_STR_RXD_LAST
--    AXI_STR_RXD_STRB
--    AXI_STR_RXD_DATA
--
--    AXI_STR_RXS_ACLK
--    AXI_STR_RXS_ARESET
--    AXI_STR_RXS_VALID
--    AXI_STR_RXS_READY
--    AXI_STR_RXS_LAST
--    AXI_STR_RXS_STRB
--    AXI_STR_RXS_DATA
--
--    EMAC_CLIENT_RXD_LEGACY
--    EMAC_CLIENT_RXD_VLD_LEGACY
--    EMAC_CLIENT_RX_GOODFRAME_LEGACY
--    EMAC_CLIENT_RX_BADFRAME_LEGACY
--    EMAC_CLIENT_RX_FRAMEDROP
--    LEGACY_RX_FILTER_MATCH
--
--    RX_CLIENT_CLK
--    RX_CLIENT_CLK_ENBL
--
--    EMAC_CLIENT_RX_STATS
--    EMAC_CLIENT_RX_STATS_VLD
--    EMAC_CLIENT_RX_STATS_BYTE_VLD
--    EMAC_CLIENT_RXD_VLD_2STATS
--    rx_statistics_vector
--
--    RTAGREGDATA
--    TPID0REGDATA
--    TPID1REGDATA
--    RX_CL_CLK_UAWL_REG_DATA
--    RX_CL_CLK_UAWU_REG_DATA
--    RXCLCLKMCASTADDR
--    RXCLCLKMCASTEN
--    RXCLCLKMCASTRDDATA
--    LLINKCLKVLANADDR
--    LLINKCLKVLANRDDATA
--    LLINKCLKRXVLANBRAMENA
--
--    LLINKCLKEMULTIFLTRENBL
--    LLINKCLKNEWFNCENBL
--    LLINKCLKRXVSTRPMODE
--    LLINKCLKRXVTAGMODE
-------------------------------------------------------------------------------
----                  Entity Section
-------------------------------------------------------------------------------

entity rx_emac_if is
    generic (
                C_RXVLAN_WIDTH        : integer                       := 12;
                C_RXD_MEM_BYTES       : integer                       := 4096;
                C_RXD_MEM_ADDR_WIDTH  : integer                       := 10;
                C_RXS_MEM_BYTES       : integer                       := 4096;
                C_RXS_MEM_ADDR_WIDTH  : integer                       := 10;
                C_ENABLE_1588          : integer   := 0;
                C_FAMILY              : string                        := "virtex6";
    C_RXCSUM              : integer range 0 to 2          := 0;
    -- 0 - No checksum offloading
    -- 1 - Partial (legacy) checksum offloading
    -- 2 - Full checksum offloading
    C_RXVLAN_TRAN         : integer range 0 to 1          := 0;
    C_RXVLAN_TAG          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP         : integer range 0 to 1          := 0;
    C_MCAST_EXTEND        : integer range 0 to 1          := 0
);

port    (
            RX_FRAME_RECEIVED_INTRPT        : out std_logic;                        --  Frame received interrupt
            RX_FRAME_REJECTED_INTRPT        : out std_logic;                        --  Frame rejected interrupt
            RX_BUFFER_MEM_OVERFLOW_INTRPT   : out std_logic;                        --  Memory overflow interrupt

            rx_statistics_vector            : in  std_logic_vector(27 downto 0);    -- RX statistics from TEMAC
            rx_statistics_valid             : in  std_logic;                        -- Rx stats valid from TEMAC
            end_of_frame_reset_in           : in  std_logic;                        -- end of frame reset base on last from rx axistream

            rx_mac_aclk                     : in  std_logic;                        -- Rx axistream clock from TEMAC
            rx_reset                        : in  std_logic;                        -- Rx axistream reset from TEMAC
            derived_rxd                     : in  std_logic_vector(7 downto 0);     -- Rx axistream data from TEMAC

            derived_rx_good_frame           : in  std_logic;                        -- derived good indicator
            derived_rx_bad_frame            : in  std_logic;                        -- derived bad indicator
            derived_rxd_vld                 : in  std_logic;                        -- derived data valid indicator
            derived_rx_clk_enbl             : in  std_logic;                        -- TEMAC clock domain enable

            RX_CL_CLK_RX_TAG_REG_DATA       : in  std_logic_vector(0 to 31);        --  Receive VLAN TAG
            RX_CL_CLK_TPID0_REG_DATA        : in  std_logic_vector(0 to 31);        --  Receive VLAN TPID 0
            RX_CL_CLK_TPID1_REG_DATA        : in  std_logic_vector(0 to 31);        --  Receive VLAN TPID 1
            RX_CL_CLK_UAWL_REG_DATA         : in  std_logic_vector(0 to 31);        --  Receive Unicast Address Word Lower
            RX_CL_CLK_UAWU_REG_DATA         : in  std_logic_vector(16 to 31);       --  Receive Unicast Address Word Upper

            RX_CL_CLK_MCAST_ADDR            : out std_logic_vector(0 to 14);        --  Receive Multicast Memory Address
            RX_CL_CLK_MCAST_EN              : out std_logic;                        --  Receive Multicast Memory Address Enable
            RX_CL_CLK_MCAST_RD_DATA         : in  std_logic_vector(0 to 0);         --  Receive Multicast Memory Address Read Data

            RX_CL_CLK_VLAN_ADDR             : out std_logic_vector(0 to 11);        --  Receive VLAN Memory Address
            RX_CL_CLK_VLAN_RD_DATA          : in  std_logic_vector(18 to 31);       --  Receive VLAN Memory Read Data
            RX_CL_CLK_VLAN_BRAM_EN_A        : out std_logic;                        --  Receive VLAN Memory Enable

            RX_CL_CLK_BAD_FRAME_ENBL        : in  std_logic;                        --  Receive Bad Frame Enable
            RX_CL_CLK_EMULTI_FLTR_ENBL      : in  std_logic;                        --  Receive Extended Multicast Address Filter Enable
            RX_CL_CLK_NEW_FNC_ENBL          : in  std_logic;                        --  Receive New Function Enable
            RX_CL_CLK_BRDCAST_REJ           : in  std_logic;                        --  Receive Broadcast Reject
            RX_CL_CLK_MULCAST_REJ           : in  std_logic;                        --  Receive Multicast Reject
            RX_CL_CLK_VSTRP_MODE            : in  std_logic_vector(0 to 1);         --  Receive VLAN Strip Mode
            RX_CL_CLK_VTAG_MODE             : in  std_logic_vector(0 to 1);         --  Receive VLAN TAG Mode

            RX_CLIENT_RXD_DPMEM_WR_DATA     : out std_logic_vector(35 downto 0);                    --  Receive Data Memory Write Data
            RX_CLIENT_RXD_DPMEM_RD_DATA     : in  std_logic_vector(35 downto 0);                    --  Receive Data Memory Read Data
            RX_CLIENT_RXD_DPMEM_WR_EN       : out std_logic_vector(0 downto 0);                     --  Receive Data Memory Write Enable
            RX_CLIENT_RXD_DPMEM_ADDR        : out std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  Receive Data Memory Address
            RX_CLIENT_RXS_DPMEM_WR_DATA     : out std_logic_vector(35 downto 0);                    --  Receive Status Memory Write Data
            RX_CLIENT_RXS_DPMEM_RD_DATA     : in  std_logic_vector(35 downto 0);                    --  Receive Status Memory Read Data
            RX_CLIENT_RXS_DPMEM_WR_EN       : out std_logic_vector(0 downto 0);                     --  Receive Status Memory Write Enable
            RX_CLIENT_RXS_DPMEM_ADDR        : out std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  Receive Status Memory Address

            AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY : in std_logic_vector(35 downto 0);    --  Receive Status Gray code pointer
            AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY : in std_logic_vector(35 downto 0)     --  Receive Data Gray code pointer
        );
end rx_emac_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of rx_emac_if is

    signal EMAC_CLIENT_RXD_LEGACY          : std_logic_vector(7 downto  0);
    signal EMAC_CLIENT_RXD_VLD_LEGACY      : std_logic;
    signal EMAC_CLIENT_RX_GOODFRAME_LEGACY : std_logic;
    signal EMAC_CLIENT_RX_BADFRAME_LEGACY  : std_logic;
    signal EMAC_CLIENT_RX_FRAMEDROP        : std_logic;
    signal LEGACY_RX_FILTER_MATCH          : std_logic_vector(7 downto 0);

    signal RX_CLIENT_CLK                   : std_logic;
    signal RX_CLIENT_CLK_ENBL              : std_logic;
    signal RESET2RX_CLIENT                 : std_logic;

    signal EMAC_CLIENT_RX_STATS            : std_logic_vector(6  downto  0);
    signal EMAC_CLIENT_RX_STATS_VLD        : std_logic;
    signal EMAC_CLIENT_RX_STATS_BYTE_VLD   : std_logic;
    signal EMAC_CLIENT_RXD_VLD_2STATS      : std_logic;
    signal SOFT_EMAC_CLIENT_RX_STATS       : std_logic_vector(27 downto 0);

---------------------------------------------------------------------
-- Functions
---------------------------------------------------------------------

-- Convert a gray code value into binary
    function gray_to_bin (
    gray : std_logic_vector)
    return std_logic_vector is

        variable binary : std_logic_vector(gray'range);

    begin

        for i in gray'high downto gray'low loop
            if i = gray'high then
                binary(i) := gray(i);
            else
                binary(i) := binary(i+1) xor gray(i);
            end if;
        end loop;  -- i

        return binary;

    end gray_to_bin;

------------------------------------------------------------------------------
-- Constant Declarations
------------------------------------------------------------------------------


------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

    type type_rx_data_words_array    is array (1 to 4) of std_logic_vector(31 downto 0);
    type type_rx_data_valid_array    is array (1 to 4) of std_logic_vector(3 downto 0);
    type type_start_of_frame_array   is array (1 to 60) of std_logic;
    type type_end_of_frame_array     is array (1 to 4) of std_logic;

    type RECEIVE_FRAME_CTRL_TYPE is (
                                    RESET_INIT_MEM_PTR_1,
                                    RESET_INIT_MEM_PTR_2,
                                    RESET_INIT_MEM_PTR_3,
                                    RESET_INIT_MEM_PTR_4,
                                    IDLE,
                                    UPDATE_MEM_PTR_1,
                                    UPDATE_STATUS_FIFO_WORD_1,
                                    UPDATE_STATUS_FIFO_WORD_2,
                                    UPDATE_STATUS_FIFO_WORD_3,
                                    UPDATE_STATUS_FIFO_WORD_4,
                                    UPDATE_STATUS_FIFO_WORD_5,
                                    UPDATE_STATUS_FIFO_WORD_6,
                                    UPDATE_MEM_PTR_2
                                );

    type RECEIVE_FRAME_DATA_TYPE is (
                                    RESET,
                                    WAIT_FOR_START_OF_FRAME,
                                    RECEIVING_FRAME,
                                    END_OF_FRAME_CHECK_GOOD_BAD
                                );


signal receive_frame_current_state : RECEIVE_FRAME_CTRL_TYPE;
signal receive_frame_next_state    : RECEIVE_FRAME_CTRL_TYPE;

signal receive_frame_data_current_state : RECEIVE_FRAME_DATA_TYPE;
signal receive_frame_data_next_state    : RECEIVE_FRAME_DATA_TYPE;

signal rx_data_words_array    : type_rx_data_words_array;
signal rx_data_valid_array    : type_rx_data_valid_array;
signal start_of_frame_array   : type_start_of_frame_array;
signal end_of_frame_array     : type_end_of_frame_array;

signal start_of_frame_d1    : std_logic;
signal save_rx_goodframe    : std_logic;
signal save_rx_badframe     : std_logic;


signal frame_is_multicast_d10           : std_logic;
signal frame_is_ip_multicast_d4         : std_logic;
signal frame_is_broadcast_d10           : std_logic;
signal first_tag_is_vlan_TPID_0_d15     : std_logic;
signal first_tag_is_vlan_TPID_1_d15     : std_logic;
signal first_tag_is_vlan_TPID_2_d15     : std_logic;
signal first_tag_is_vlan_TPID_3_d15     : std_logic;
signal second_tag_is_vlan_TPID_0_d19    : std_logic;
signal second_tag_is_vlan_TPID_1_d19    : std_logic;
signal second_tag_is_vlan_TPID_2_d19    : std_logic;
signal second_tag_is_vlan_TPID_3_d19    : std_logic;
signal frame_is_vlan_8100_d15           : std_logic;
signal frame_has_valid_length_field_d22 : std_logic;
signal frame_has_type_0800_d22          : std_logic;
signal frame_is_snap_d30                : std_logic;
signal frame_is_ip_protocol_d31         : std_logic;
signal frame_has_ip_hdr_length_d31      : std_logic;
signal frame_has_no_ip_frags_d38        : std_logic;
signal frame_has_udp_protocol_d38       : std_logic;
signal frame_has_tcp_protocol_d38       : std_logic;
signal pack_high_1_pack_low_0           : std_logic;
signal rxd_packed_16bits                : unsigned(15 downto 0);
signal enable_ip_hdr_sum_1              : std_logic;
signal ip_header_sum_1                  : unsigned(16 downto 0);
signal enable_ip_hdr_sum_2              : std_logic;
signal ip_header_sum_2                  : unsigned(16 downto 0);
signal enable_ip_hdr_sum_3              : std_logic;
signal ip_header_sum_3                  : unsigned(16 downto 0);
signal enable_ip_hdr_sum_4              : std_logic;
signal ip_header_sum_4                  : unsigned(16 downto 0);
signal ip_header_csum_1_ok              : std_logic;
signal ip_header_csum_2_ok              : std_logic;
signal ip_header_csum_3_ok              : std_logic;
signal ip_header_csum_4_ok              : std_logic;
signal frame_ip_csum_checked            : std_logic;
signal frame_udp_csum_checked           : std_logic;
signal frame_tcp_csum_checked           : std_logic;
signal frame_is_e2                      : std_logic;
signal frame_is_e2_vlan                 : std_logic;
signal frame_is_snap                    : std_logic;
signal frame_is_snap_vlan               : std_logic;
signal frame_ip_csum_ok                 : std_logic;
signal frame_udp_csum_ok                : std_logic;
signal frame_tcp_csum_ok                : std_logic;
signal receive_checksum_status          : std_logic_vector(2 downto 0);
signal receive_checksum_status_i        : std_logic_vector(2 downto 0);

signal enable_udp_hdr_sum_1             : std_logic;
signal udp_header_sum_1                 : unsigned(16 downto 0);
signal udp_header_csum_1_ok             : std_logic;
signal save_udp_hdr_length_1            : std_logic_vector(15 downto 0);
signal enable_udp_hdr_sum_2             : std_logic;
signal udp_header_sum_2                 : unsigned(16 downto 0);
signal udp_header_csum_2_ok             : std_logic;
signal save_udp_hdr_length_2            : std_logic_vector(15 downto 0);
signal enable_udp_hdr_sum_3             : std_logic;
signal udp_header_sum_3                 : unsigned(16 downto 0);
signal udp_header_csum_3_ok             : std_logic;
signal save_udp_hdr_length_3            : std_logic_vector(15 downto 0);
signal enable_udp_hdr_sum_4             : std_logic;
signal udp_header_sum_4                 : unsigned(16 downto 0);
signal udp_header_csum_4_ok             : std_logic;
signal save_udp_hdr_length_4            : std_logic_vector(15 downto 0);

signal save_tcp_length_1                : std_logic_vector(15 downto 0);
signal enable_tcp_hdr_sum_1             : std_logic;
signal tcp_header_sum_1                 : unsigned(16 downto 0);
signal tcp_header_csum_1_ok             : std_logic;
signal save_tcp_length_2                : std_logic_vector(15 downto 0);
signal enable_tcp_hdr_sum_2             : std_logic;
signal tcp_header_sum_2                 : unsigned(16 downto 0);
signal tcp_header_csum_2_ok             : std_logic;
signal save_tcp_length_3                : std_logic_vector(15 downto 0);
signal enable_tcp_hdr_sum_3             : std_logic;
signal tcp_header_sum_3                 : unsigned(16 downto 0);
signal tcp_header_csum_3_ok             : std_logic;
signal save_tcp_length_4                : std_logic_vector(15 downto 0);
signal enable_tcp_hdr_sum_4             : std_logic;
signal tcp_header_sum_4                 : unsigned(16 downto 0);
signal tcp_header_csum_4_ok             : std_logic;

signal rx_data_packed_word              : std_logic_vector(31 downto 0);
signal rx_data_vld_packed_word          : std_logic_vector(3 downto 0);
signal rx_data_packed_state             : std_logic_vector(1 downto 0);
signal rx_data_packed_ready             : std_logic;

signal frame_length_bytes               : unsigned(15 downto 0);
signal frame_length_bytes_lat           : unsigned(15 downto 0);

signal rxd_mem_next_available4write_ptr_cmb : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_next_available4write_ptr_reg : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_last_read_out_ptr_cmb        : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_last_read_out_ptr_reg        : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_next_available4write_ptr_cmb : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_next_available4write_ptr_reg : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);

signal rxd_mem_full_mask                : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_full_mask_minus_one      : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_empty_mask               : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_one_mask                 : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_two_mask                 : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_full_mask                : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_full_mask_minus_one      : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_empty_mask               : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_one_mask                 : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_two_mask                 : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_three_mask               : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_four_mask                : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);

signal zero_extend_rxd_mask36           : std_logic_vector(35 downto C_RXD_MEM_ADDR_WIDTH + 1);
signal zero_extend_rxs_mask36           : std_logic_vector(35 downto C_RXS_MEM_ADDR_WIDTH + 1);

signal rxs_status_word_1_cmb            : std_logic_vector(35 downto 0);
signal rxs_status_word_1_reg            : std_logic_vector(35 downto 0);
signal rxs_status_word_2                : std_logic_vector(35 downto 0);
signal rxs_status_word_3                : std_logic_vector(35 downto 0);
signal rxs_status_word_4                : std_logic_vector(35 downto 0);
signal rxs_status_word_5                : std_logic_vector(35 downto 0);
signal rxs_status_word_6_cmb            : std_logic_vector(35 downto 0);
signal rxs_status_word_6_reg            : std_logic_vector(35 downto 0);

signal rxd_addr_cntr_en                 : std_logic;
signal rxs_addr_cntr_en                 : std_logic;
signal rxd_mem_addr_cntr                : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_addr_cntr                : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxd_addr_cntr_load               : std_logic;
signal rxs_addr_cntr_load               : std_logic;
signal update_status_fifo               : std_logic;

signal multicast_addr_upper_d10         : std_logic_vector(15 downto 0);
signal multicast_addr_lower_d10         : std_logic_vector(31 downto 0);
signal bytes_12_and_13_d19              : std_logic_vector(15 downto 0);
signal bytes_14_and_15_d19              : std_logic_vector(15 downto 0);

signal raw_checksum                     : std_logic_vector(15 downto 0);

signal statistics_vector                : std_logic_vector(25 downto 0);
signal frame_drop                       : std_logic;
signal not_enough_rxs_memory            : std_logic;

signal rxCsum                           : std_logic_vector(15 downto 0);
signal rxCsumVld                        : std_logic;


signal extendedMulticastReject          : std_logic;
signal saveExtendedMulticastReject : std_logic;

signal rxclclk_rxd_mem_last_read_out_ptr           : std_logic_vector(35 downto 0);
signal rxclclk_rxd_mem_last_read_out_ptr_d1        : std_logic_vector(35 downto 0);
signal sync_rxd_mem_last_read_out_ptr_gray_sync    : std_logic_vector(35 downto 0);

signal rxclclk_rxs_mem_last_read_out_ptr           : unsigned(35 downto 0);
signal rxclclk_rxs_mem_last_read_out_ptr_d1        : unsigned(35 downto 0);
signal sync_rxs_mem_last_read_out_ptr_gray_sync    : std_logic_vector(35 downto 0);

signal eof_reset : std_logic;

signal udp_pack_len_cntr_1 : unsigned(15 downto 0);
signal udp_len_is_odd_1    : std_logic;
signal udp_eof_reached_1   : std_logic;
signal udp_pack_len_cntr_2 : unsigned(15 downto 0);
signal udp_len_is_odd_2    : std_logic;
signal udp_eof_reached_2   : std_logic;
signal udp_pack_len_cntr_3 : unsigned(15 downto 0);
signal udp_len_is_odd_3    : std_logic;
signal udp_eof_reached_3   : std_logic;
signal udp_pack_len_cntr_4 : unsigned(15 downto 0);
signal udp_len_is_odd_4    : std_logic;
signal udp_eof_reached_4   : std_logic;

signal tcp_pack_len_cntr_1 : unsigned(15 downto 0);
signal tcp_len_is_odd_1    : std_logic;
signal tcp_eof_reached_1   : std_logic;
signal tcp_pack_len_cntr_2 : unsigned(15 downto 0);
signal tcp_len_is_odd_2    : std_logic;
signal tcp_eof_reached_2   : std_logic;
signal tcp_pack_len_cntr_3 : unsigned(15 downto 0);
signal tcp_len_is_odd_3    : std_logic;
signal tcp_eof_reached_3   : std_logic;
signal tcp_pack_len_cntr_4 : unsigned(15 downto 0);
signal tcp_len_is_odd_4    : std_logic;
signal tcp_eof_reached_4   : std_logic;
signal initial_index       : integer;


begin

    EMAC_CLIENT_RXD_VLD_LEGACY      <= derived_rxd_vld;
    RX_CLIENT_CLK_ENBL              <= derived_rx_clk_enbl;

    EMAC_CLIENT_RX_GOODFRAME_LEGACY <= derived_rx_good_frame;
    EMAC_CLIENT_RX_BADFRAME_LEGACY  <= derived_rx_bad_frame;
    EMAC_CLIENT_RX_STATS_VLD        <= rx_statistics_valid;
    SOFT_EMAC_CLIENT_RX_STATS       <= rx_statistics_vector;
    RX_CLIENT_CLK                   <= rx_mac_aclk;
    RESET2RX_CLIENT                 <= rx_reset;
    EMAC_CLIENT_RXD_LEGACY          <= derived_rxd;

    eof_reset <= end_of_frame_reset_in;

    ENABLE_ZERO_INIT_CNT: if(C_ENABLE_1588 = 0) generate
    begin 
	initial_index <= 0;
    end generate ENABLE_ZERO_INIT_CNT;

    ENABLE_EIGHT_INIT_CNT: if(C_ENABLE_1588 > 0) generate
    begin 
	initial_index <= 8;
    end generate ENABLE_EIGHT_INIT_CNT;

    NO_FULL_CSUM_OFFLOAD: if(not(C_RXCSUM = 2)) generate
    begin
        receive_checksum_status  <= "000";
    end generate NO_FULL_CSUM_OFFLOAD;

    YES_FULL_CSUM_OFFLOAD: if (C_RXCSUM = 2) generate
    begin
        receive_checksum_status_i <= "000" when frame_ip_csum_checked  = '0' else
                                     "001" when frame_ip_csum_checked  = '1' and frame_ip_csum_ok = '1' and frame_udp_csum_checked = '0' and frame_tcp_csum_checked = '0' else
                                     "010" when frame_ip_csum_checked  = '1' and frame_ip_csum_ok = '1' and frame_tcp_csum_checked = '1' and frame_tcp_csum_ok = '1' else
                                     "011" when frame_ip_csum_checked  = '1' and frame_ip_csum_ok = '1' and frame_udp_csum_checked = '1' and frame_udp_csum_ok = '1' else
                                     "101" when frame_ip_csum_checked  = '1' and frame_ip_csum_ok = '0' else
                                     "110" when frame_ip_csum_checked  = '1' and frame_ip_csum_ok = '1' and frame_tcp_csum_checked = '1' and frame_tcp_csum_ok = '0' else
                                     "111" when frame_ip_csum_checked  = '1' and frame_ip_csum_ok = '1' and frame_udp_csum_checked = '1' and frame_udp_csum_ok = '0' else
                                     "100"; -- should never get this value!

        REG_CSUM_STATUS_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    receive_checksum_status  <= "000";
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            receive_checksum_status  <= "000";
                        else
                            receive_checksum_status  <= receive_checksum_status_i;
                        end if;
                    end if;
                end if;
            end if;
        end process;

        IP_CSUM_CHECKED_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_ip_csum_checked  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_ip_csum_checked  <= '0';
                        elsif (frame_has_type_0800_d22 = '1' or frame_is_snap_d30 = '1') and frame_has_ip_hdr_length_d31 = '1' and
                        frame_is_ip_protocol_d31 = '1' and frame_has_no_ip_frags_d38 = '1' then
                            frame_ip_csum_checked  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        UDP_CSUM_CHECKED_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_udp_csum_checked  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_udp_csum_checked  <= '0';
                        elsif frame_ip_csum_checked = '1' and frame_has_udp_protocol_d38 = '1' and frame_ip_csum_checked = '1' and
                        frame_ip_csum_ok = '1' then
                            frame_udp_csum_checked  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        TCP_CSUM_CHECKED_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_tcp_csum_checked  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_tcp_csum_checked  <= '0';
                        elsif frame_ip_csum_checked = '1' and frame_has_tcp_protocol_d38 = '1' and frame_ip_csum_checked = '1' and frame_ip_csum_ok = '1' then
                            frame_tcp_csum_checked  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        FRAME_IS_ETHERNET_2_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_is_e2  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_is_e2  <= '0';
                        elsif frame_has_type_0800_d22 = '1' and frame_is_vlan_8100_d15 = '0' then
                            frame_is_e2  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        FRAME_IS_ETHERNET_2VLAN_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_is_e2_vlan  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_is_e2_vlan  <= '0';
                        elsif frame_has_type_0800_d22 = '1' and frame_is_vlan_8100_d15 = '1' then
                            frame_is_e2_vlan  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        FRAME_IS_SNAP_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_is_snap  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_is_snap  <= '0';
                        elsif frame_is_snap_d30 = '1' and frame_is_vlan_8100_d15 = '0' then
                            frame_is_snap  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        FRAME_IS_SNAPVLAN_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_is_snap_vlan  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_is_snap_vlan  <= '0';
                        elsif frame_is_snap_d30 = '1' and frame_is_vlan_8100_d15 = '1' then
                            frame_is_snap_vlan  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        IP_CSUM_IS_OK_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_ip_csum_ok  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_ip_csum_ok  <= '0';
                        elsif frame_ip_csum_checked = '1' and ((frame_is_e2 = '1'        and ip_header_csum_1_ok = '1') or
                        (frame_is_e2_vlan = '1'   and ip_header_csum_2_ok = '1') or
                        (frame_is_snap = '1'      and ip_header_csum_3_ok = '1') or
                        (frame_is_snap_vlan = '1' and ip_header_csum_4_ok = '1')) then
                            frame_ip_csum_ok  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        UDP_CSUM_IS_OK_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_udp_csum_ok  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_udp_csum_ok  <= '0';
                        elsif frame_udp_csum_checked = '1' and 
                            ((frame_is_e2 = '1'       and udp_header_csum_1_ok = '1') or
                            (frame_is_e2_vlan = '1'   and udp_header_csum_2_ok = '1') or
                            (frame_is_snap = '1'      and udp_header_csum_3_ok = '1') or
                            (frame_is_snap_vlan = '1' and udp_header_csum_4_ok = '1')) then
                            frame_udp_csum_ok  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        TCP_CSUM_IS_OK_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_tcp_csum_ok  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if(eof_reset = '1') then
                            frame_tcp_csum_ok  <= '0';
                        elsif frame_tcp_csum_checked = '1' and ((frame_is_e2 = '1'        and tcp_header_csum_1_ok = '1') or
                        (frame_is_e2_vlan = '1'   and tcp_header_csum_2_ok = '1') or
                        (frame_is_snap = '1'      and tcp_header_csum_3_ok = '1') or
                        (frame_is_snap_vlan = '1' and tcp_header_csum_4_ok = '1')) then
                            frame_tcp_csum_ok  <= '1';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_IP_HDR_1_PROCESS: process (RX_CLIENT_CLK) -- no vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    ip_header_sum_1  <=(others => '0');
                    ip_header_csum_1_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            ip_header_csum_1_ok <= '0';
                        elsif (ip_header_sum_1(15 downto 0) = X"FFFF" and ip_header_sum_1(16) = '0' and enable_ip_hdr_sum_1 = '0') then
                            ip_header_csum_1_ok <= '1';
                        else
                            ip_header_csum_1_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            ip_header_sum_1  <=(others => '0');
                        elsif (enable_ip_hdr_sum_1 = '1' and pack_high_1_pack_low_0 = '1') then
                            ip_header_sum_1(16 downto 0)  <= ('0'&ip_header_sum_1(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                        elsif (enable_ip_hdr_sum_1 = '1' and pack_high_1_pack_low_0 = '0') then
                            -- wrap previous carry back in
                            ip_header_sum_1(16 downto 0)  <= ('0'&ip_header_sum_1(15 downto 0)) + (X"0000"&ip_header_sum_1(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        ENABLE_IP_HEADER_SUM_1_PROCESS: process (RX_CLIENT_CLK) -- no vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_ip_hdr_sum_1  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 15) = '1') then
                            enable_ip_hdr_sum_1  <= '1';
                        elsif(start_of_frame_array(initial_index + 35) = '1') then
                            enable_ip_hdr_sum_1  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_IP_HDR_2_PROCESS: process (RX_CLIENT_CLK) -- yes vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    ip_header_sum_2  <=(others => '0');
                    ip_header_csum_2_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            ip_header_csum_2_ok <= '0';
                        elsif (ip_header_sum_2(15 downto 0) = X"FFFF" and ip_header_sum_2(16) = '0' and enable_ip_hdr_sum_2 = '0') then
                            ip_header_csum_2_ok <= '1';
                        else
                            ip_header_csum_2_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            ip_header_sum_2  <=(others => '0');
                        elsif (enable_ip_hdr_sum_2 = '1' and pack_high_1_pack_low_0 = '1') then
                            ip_header_sum_2(16 downto 0)  <= ('0'&ip_header_sum_2(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                        elsif (enable_ip_hdr_sum_2 = '1' and pack_high_1_pack_low_0 = '0') then
                            -- wrap previous carry back in
                            ip_header_sum_2(16 downto 0)  <= ('0'&ip_header_sum_2(15 downto 0)) + (X"0000"&ip_header_sum_2(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        ENABLE_IP_HEADER_SUM_2_PROCESS: process (RX_CLIENT_CLK) -- yes vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_ip_hdr_sum_2 <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 19) = '1') then
                            enable_ip_hdr_sum_2  <= '1';
                        elsif(start_of_frame_array(initial_index + 39) = '1') then
                            enable_ip_hdr_sum_2  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_IP_HDR_3_PROCESS: process (RX_CLIENT_CLK) -- no vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    ip_header_sum_3  <=(others => '0');
                    ip_header_csum_3_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            ip_header_csum_3_ok <= '0';
                        elsif (ip_header_sum_3(15 downto 0) = X"FFFF" and ip_header_sum_3(16) = '0' and enable_ip_hdr_sum_3 = '0') then
                            ip_header_csum_3_ok <= '1';
                        else
                            ip_header_csum_3_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            ip_header_sum_3  <=(others => '0');
                        elsif (enable_ip_hdr_sum_3 = '1' and pack_high_1_pack_low_0 = '1') then
                            ip_header_sum_3(16 downto 0)  <= ('0'&ip_header_sum_3(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                        elsif (enable_ip_hdr_sum_3 = '1' and pack_high_1_pack_low_0 = '0') then
                            -- wrap previous carry back in
                            ip_header_sum_3(16 downto 0)  <= ('0'&ip_header_sum_3(15 downto 0)) + (X"0000"&ip_header_sum_3(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        ENABLE_IP_HEADER_SUM_3_PROCESS: process (RX_CLIENT_CLK) -- no vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_ip_hdr_sum_3  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 23) = '1') then
                            enable_ip_hdr_sum_3  <= '1';
                        elsif(start_of_frame_array(initial_index + 43) = '1') then
                            enable_ip_hdr_sum_3  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_IP_HDR_4_PROCESS: process (RX_CLIENT_CLK) -- yes vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    ip_header_sum_4  <=(others => '0');
                    ip_header_csum_4_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            ip_header_csum_4_ok <= '0';
                        elsif (ip_header_sum_4(15 downto 0) = X"FFFF" and ip_header_sum_4(16) = '0' and enable_ip_hdr_sum_4 = '0') then
                            ip_header_csum_4_ok <= '1';
                        else
                            ip_header_csum_4_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            ip_header_sum_4  <=(others => '0');
                        elsif (enable_ip_hdr_sum_4 = '1' and pack_high_1_pack_low_0 = '1') then
                            ip_header_sum_4(16 downto 0)  <= ('0'&ip_header_sum_4(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                        elsif (enable_ip_hdr_sum_4 = '1' and pack_high_1_pack_low_0 = '0') then
                            -- wrap previous carry back in
                            ip_header_sum_4(16 downto 0)  <= ('0'&ip_header_sum_4(15 downto 0)) + (X"0000"&ip_header_sum_4(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        ENABLE_IP_HEADER_SUM_4_PROCESS: process (RX_CLIENT_CLK) -- yes vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_ip_hdr_sum_4  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 27) = '1') then
                            enable_ip_hdr_sum_4  <= '1';
                        elsif(start_of_frame_array(initial_index + 47) = '1') then
                            enable_ip_hdr_sum_4  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_UDP_HDR_1_PROCESS: process (RX_CLIENT_CLK) -- no vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    udp_header_sum_1  <=(others => '0');
                    udp_header_csum_1_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            udp_header_csum_1_ok <= '0';
                        elsif ((udp_header_sum_1(15 downto 0) + unsigned(save_udp_hdr_length_1)) = X"FFFF" and udp_header_sum_1(16) = '0' and enable_udp_hdr_sum_1 = '0') then
                            udp_header_csum_1_ok <= '1';
                        elsif ((udp_header_sum_1(15 downto 0) + unsigned(save_udp_hdr_length_1)) = X"FFFE" and udp_header_sum_1(16) = '1' and enable_udp_hdr_sum_1 = '0') then
                            udp_header_csum_1_ok <= '1';
                        else
                            udp_header_csum_1_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            udp_header_sum_1  <=(others => '0');
                        elsif (enable_udp_hdr_sum_1 = '1' and pack_high_1_pack_low_0 = '1') then
                            if (start_of_frame_array(initial_index + 24) = '1') then -- mask Time to live filed from protocol in Ip header
                                udp_header_sum_1(16 downto 0)  <= ('0'&udp_header_sum_1(15 downto 0)) + ("000000000"&rxd_packed_16bits(7 downto 0));
                            elsif (start_of_frame_array(initial_index + 26) = '1') then -- mask IP header csum
                                udp_header_sum_1(16 downto 0)  <= ('0'&udp_header_sum_1(15 downto 0));
                            elsif(udp_eof_reached_1 = '1' and udp_len_is_odd_1 = '1') then
              -- In case of Odd-length UDP packet, for last checksum word input, the LSB is padded with Zeros
                                udp_header_sum_1(16 downto 0)  <= ('0' & udp_header_sum_1(15 downto 0)) + (rxd_packed_16bits(15 downto 8) & x"00");
                            else
                                udp_header_sum_1(16 downto 0)  <= ('0'&udp_header_sum_1(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                            end if;
                        elsif (enable_udp_hdr_sum_1 = '1' and pack_high_1_pack_low_0 = '0') then
            -- wrap previous carry back in
                            udp_header_sum_1(16 downto 0)  <= ('0'&udp_header_sum_1(15 downto 0)) + (X"0000"&udp_header_sum_1(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SAVE_UDP_HEADER_LENGTH_1_PROCESS: process (RX_CLIENT_CLK) -- no vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    save_udp_hdr_length_1  <= (others => '0');
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 40) = '1') then
                            save_udp_hdr_length_1  <= std_logic_vector(rxd_packed_16bits);
                        elsif(eof_reset = '1') then
                            save_udp_hdr_length_1  <= (others => '0');
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -- Counter to track the #2-byte words from UDP packet to be used for checksum calculation
        udp_pack_len_cntr_1_process: process(rx_client_clk)
            variable udp_pack_len_cntr_1_div2 : unsigned(15 downto 0);
        begin
            if(rising_edge(rx_client_clk)) then
                if(reset2rx_client = '1' or eof_reset = '1') then
                    udp_pack_len_cntr_1 <= (others => '1');
                elsif(rx_client_clk_enbl = '1' and start_of_frame_array(initial_index + 40) = '1') then
          -- Load the counter with the UDP packet length and discount the #2-byte words till this point in time
          -- Counter Value = (UDP Pack Len/2) - 3. (#2-byte words already added to Checksum Calculation)
                    udp_pack_len_cntr_1_div2  := '0' & rxd_packed_16bits(15 downto 1);
                    udp_pack_len_cntr_1       <= udp_pack_len_cntr_1_div2-x"0003";   
                elsif(rx_client_clk_enbl = '1' and udp_pack_len_cntr_1 /= x"FFFF" and enable_udp_hdr_sum_1 = '1' and pack_high_1_pack_low_0 = '1') then
                    udp_pack_len_cntr_1 <= udp_pack_len_cntr_1-x"0001";
                end if;
            end if;
        end process;

        udp_len_is_odd_1  <= save_udp_hdr_length_1(0);
        udp_eof_reached_1 <= '1' when ((udp_pack_len_cntr_1 = x"0001" and udp_len_is_odd_1 = '0') or (udp_pack_len_cntr_1 = x"0000" and udp_len_is_odd_1 = '1')) 
                             else '0'; 

        ENABLE_UDP_HEADER_SUM_1_PROCESS: process (RX_CLIENT_CLK) -- no vlan no snap 
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_udp_hdr_sum_1  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 23) = '1') then
                            enable_udp_hdr_sum_1  <= '1';
                        elsif((udp_eof_reached_1 = '1' and pack_high_1_pack_low_0 = '1') or start_of_frame_d1 = '0') then
                            enable_udp_hdr_sum_1  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_UDP_HDR_2_PROCESS: process (RX_CLIENT_CLK) -- yes vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    udp_header_sum_2  <=(others => '0');
                    udp_header_csum_2_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            udp_header_csum_2_ok <= '0';
                        elsif ((udp_header_sum_2(15 downto 0) + unsigned(save_udp_hdr_length_2)) = X"FFFF" and udp_header_sum_2(16) = '0' and
                        enable_udp_hdr_sum_2 = '0') then
                            udp_header_csum_2_ok <= '1';
                        elsif ((udp_header_sum_2(15 downto 0) + unsigned(save_udp_hdr_length_2)) = X"FFFE" and udp_header_sum_2(16) = '1' and
                        enable_udp_hdr_sum_2 = '0') then
                            udp_header_csum_2_ok <= '1';
                        else
                            udp_header_csum_2_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            udp_header_sum_2  <=(others => '0');
                        elsif (enable_udp_hdr_sum_2 = '1' and pack_high_1_pack_low_0 = '1') then
                            if (start_of_frame_array(initial_index + 28) = '1') then -- mask Time to live filed from protocol in Ip header
                                udp_header_sum_2(16 downto 0)  <= ('0'&udp_header_sum_2(15 downto 0)) + ("000000000"&rxd_packed_16bits(7 downto 0));
                            elsif (start_of_frame_array(initial_index + 30) = '1') then -- mask IP header csum
                                udp_header_sum_2(16 downto 0)  <= ('0'&udp_header_sum_2(15 downto 0)) + ("00000000000000000");
                            elsif(udp_eof_reached_2 = '1' and udp_len_is_odd_2 = '1') then
              -- In case of Odd-length UDP packet, for last checksum word input, the LSB is padded with Zeros
                                udp_header_sum_2(16 downto 0)  <= ('0'&udp_header_sum_2(15 downto 0)) + (rxd_packed_16bits(15 downto 8) & x"00");
                            else
                                udp_header_sum_2(16 downto 0)  <= ('0'&udp_header_sum_2(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                            end if;
                        elsif (enable_udp_hdr_sum_2 = '1' and pack_high_1_pack_low_0 = '0') then
            -- wrap previous carry back in
                            udp_header_sum_2(16 downto 0)  <= ('0'&udp_header_sum_2(15 downto 0)) + (X"0000"&udp_header_sum_2(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SAVE_UDP_HEADER_LENGTH_2_PROCESS: process (RX_CLIENT_CLK) -- yes vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    save_udp_hdr_length_2  <= (others => '0');
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 44) = '1') then
                            save_udp_hdr_length_2  <= std_logic_vector(rxd_packed_16bits);
                        elsif(eof_reset = '1') then
                            save_udp_hdr_length_2  <= (others => '0');
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -- Counter to track the #2-byte words from UDP packet to be used for checksum calculation
        udp_pack_len_cntr_2_process: process(rx_client_clk)
            variable udp_pack_len_cntr_2_div2 : unsigned(15 downto 0);
        begin
            if(rising_edge(rx_client_clk)) then
                if(reset2rx_client = '1' or eof_reset = '1') then
                    udp_pack_len_cntr_2 <= (others => '0');
                elsif(rx_client_clk_enbl = '1' and start_of_frame_array(initial_index + 44) = '1') then
          -- Load the counter with the UDP packet length and discount the #2-byte words till this point in time
          -- Counter Value = (UDP Pack Len/2) - 3. (#2-byte words already added to Checksum Calculation)
                    udp_pack_len_cntr_2_div2  := '0' & rxd_packed_16bits(15 downto 1);
                    udp_pack_len_cntr_2       <= udp_pack_len_cntr_2_div2-x"0003";   
                elsif(rx_client_clk_enbl = '1' and udp_pack_len_cntr_2 /= x"FFFF" and enable_udp_hdr_sum_2 = '1' and pack_high_1_pack_low_0 = '1') then
                    udp_pack_len_cntr_2 <= udp_pack_len_cntr_2-x"0001";
                end if;
            end if;
        end process;

        udp_len_is_odd_2  <= save_udp_hdr_length_2(0);
        udp_eof_reached_2 <= '1' when ((udp_pack_len_cntr_2 = x"0001" and udp_len_is_odd_2 = '0') or (udp_pack_len_cntr_2 = x"0000" and udp_len_is_odd_2= '1')) 
                             else '0'; 

        ENABLE_UDP_HEADER_SUM_2_PROCESS: process (RX_CLIENT_CLK) -- yes vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_udp_hdr_sum_2  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 27) = '1') then
                            enable_udp_hdr_sum_2  <= '1';
                        elsif((udp_eof_reached_2 = '1' and pack_high_1_pack_low_0 = '1') or start_of_frame_d1 = '0') then
                            enable_udp_hdr_sum_2  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_UDP_HDR_3_PROCESS: process (RX_CLIENT_CLK) -- no vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    udp_header_sum_3  <=(others => '0');
                    udp_header_csum_3_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            udp_header_csum_3_ok <= '0';
                        elsif ((udp_header_sum_3(15 downto 0) + unsigned(save_udp_hdr_length_3)) = X"FFFF" and udp_header_sum_3(16) = '0' and
                        enable_udp_hdr_sum_3 = '0') then
                            udp_header_csum_3_ok <= '1';
                        elsif ((udp_header_sum_3(15 downto 0) + unsigned(save_udp_hdr_length_3)) = X"FFFE" and udp_header_sum_3(16) = '1' and
                        enable_udp_hdr_sum_3 = '0') then
                            udp_header_csum_3_ok <= '1';
                        else
                            udp_header_csum_3_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            udp_header_sum_3  <=(others => '0');
                        elsif (enable_udp_hdr_sum_3 = '1' and pack_high_1_pack_low_0 = '1') then
                            if (start_of_frame_array(initial_index + 32) = '1') then -- mask Time to live filed from protocol in Ip header
                                udp_header_sum_3(16 downto 0)  <= ('0'&udp_header_sum_3(15 downto 0)) + ("000000000"&rxd_packed_16bits(7 downto 0));
                            elsif (start_of_frame_array(initial_index + 34) = '1') then -- mask IP header csum
                                udp_header_sum_3(16 downto 0)  <= ('0'&udp_header_sum_3(15 downto 0)) + ("00000000000000000");
                            elsif(udp_eof_reached_3 = '1' and udp_len_is_odd_3 = '1') then
              -- In case of Odd-length UDP packet, for last checksum word input, the LSB is padded with Zeros
                                udp_header_sum_3(16 downto 0)  <= ('0'&udp_header_sum_3(15 downto 0)) + (rxd_packed_16bits(15 downto 8) & x"00");
                            else
                                udp_header_sum_3(16 downto 0)  <= ('0'&udp_header_sum_3(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                            end if;
                        elsif (enable_udp_hdr_sum_3 = '1' and pack_high_1_pack_low_0 = '0') then
            -- wrap previous carry back in
                            udp_header_sum_3(16 downto 0)  <= ('0'&udp_header_sum_3(15 downto 0)) + (X"0000"&udp_header_sum_3(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SAVE_UDP_HEADER_LENGTH_3_PROCESS: process (RX_CLIENT_CLK) -- no vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    save_udp_hdr_length_3  <= (others => '0');
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 48) = '1') then
                            save_udp_hdr_length_3  <= std_logic_vector(rxd_packed_16bits);
                        elsif(eof_reset = '1') then
                            save_udp_hdr_length_3  <= (others => '0');
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -- Counter to track the #2-byte words from UDP packet to be used for checksum calculation
        udp_pack_len_cntr_3_process: process(rx_client_clk)
            variable udp_pack_len_cntr_3_div2 : unsigned(15 downto 0);
        begin
            if(rising_edge(rx_client_clk)) then
                if(reset2rx_client = '1' or eof_reset = '1') then
                    udp_pack_len_cntr_3 <= (others => '1');
                elsif(rx_client_clk_enbl = '1' and start_of_frame_array(initial_index + 48) = '1') then
          -- Load the counter with the UDP packet length and discount the #2-byte words till this point in time
          -- Counter Value = (UDP Pack Len/2) - 3. (#2-byte words already added to Checksum Calculation)
                    udp_pack_len_cntr_3_div2  := '0' & rxd_packed_16bits(15 downto 1);
                    udp_pack_len_cntr_3       <= udp_pack_len_cntr_3_div2-x"0003";   
                elsif(rx_client_clk_enbl = '1' and udp_pack_len_cntr_3 /= x"FFFF" and enable_udp_hdr_sum_3 = '1' and pack_high_1_pack_low_0 = '1') then
                    udp_pack_len_cntr_3 <= udp_pack_len_cntr_3-x"0001";
                end if;
            end if;
        end process;

        udp_len_is_odd_3  <= save_udp_hdr_length_3(0);
        udp_eof_reached_3 <= '1' when ((udp_pack_len_cntr_3 = x"0001" and udp_len_is_odd_3 = '0') or (udp_pack_len_cntr_3 = x"0000" and udp_len_is_odd_3 = '1')) 
                             else '0'; 

        ENABLE_UDP_HEADER_SUM_3_PROCESS: process (RX_CLIENT_CLK) -- no vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_udp_hdr_sum_3  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 31) = '1') then
                            enable_udp_hdr_sum_3  <= '1';
                        elsif((udp_eof_reached_3 = '1' and pack_high_1_pack_low_0 = '1') or start_of_frame_d1 = '0') then
                            enable_udp_hdr_sum_3  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_UDP_HDR_4_PROCESS: process (RX_CLIENT_CLK) -- yes vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    udp_header_sum_4  <=(others => '0');
                    udp_header_csum_4_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            udp_header_csum_4_ok <= '0';
                        elsif ((udp_header_sum_4(15 downto 0) + unsigned(save_udp_hdr_length_4)) = X"FFFF" and udp_header_sum_4(16) = '0' and
                        enable_udp_hdr_sum_4 = '0') then
                            udp_header_csum_4_ok <= '1';
                        elsif ((udp_header_sum_4(15 downto 0) + unsigned(save_udp_hdr_length_4)) = X"FFFE" and udp_header_sum_4(16) = '1' and
                        enable_udp_hdr_sum_4 = '0') then
                            udp_header_csum_4_ok <= '1';
                        else
                            udp_header_csum_4_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            udp_header_sum_4  <=(others => '0');
                        elsif (enable_udp_hdr_sum_4 = '1' and pack_high_1_pack_low_0 = '1') then
                            if (start_of_frame_array(initial_index + 36) = '1') then -- mask Time to live filed from protocol in Ip header
                                udp_header_sum_4(16 downto 0)  <= ('0'&udp_header_sum_4(15 downto 0)) + ("000000000"&rxd_packed_16bits(7 downto 0));
                            elsif (start_of_frame_array(initial_index + 38) = '1') then -- mask IP header csum
                                udp_header_sum_4(16 downto 0)  <= ('0'&udp_header_sum_4(15 downto 0)) + ("00000000000000000");
                            elsif(udp_eof_reached_4 = '1' and udp_len_is_odd_4 = '1') then
              -- In case of Odd-length UDP packet, for last checksum word input, the LSB is padded with Zeros
                                udp_header_sum_4(16 downto 0)  <= ('0'&udp_header_sum_4(15 downto 0)) + (rxd_packed_16bits(15 downto 8) & x"00");
                            else
                                udp_header_sum_4(16 downto 0)  <= ('0'&udp_header_sum_4(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                            end if;
                        elsif (enable_udp_hdr_sum_4 = '1' and pack_high_1_pack_low_0 = '0') then
            -- wrap previous carry back in
                            udp_header_sum_4(16 downto 0)  <= ('0'&udp_header_sum_4(15 downto 0)) + (X"0000"&udp_header_sum_4(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SAVE_UDP_HEADER_LENGTH_4_PROCESS: process (RX_CLIENT_CLK) -- yes vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    save_udp_hdr_length_4  <= (others => '0');
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 52) = '1') then
                            save_udp_hdr_length_4  <= std_logic_vector(rxd_packed_16bits);
                        elsif(eof_reset = '1') then
                            save_udp_hdr_length_4  <= (others => '0');
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -- Counter to track the #2-byte words from UDP packet to be used for checksum calculation
        udp_pack_len_cntr_4_process: process(rx_client_clk)
            variable udp_pack_len_cntr_4_div2 : unsigned(15 downto 0);
        begin
            if(rising_edge(rx_client_clk)) then
                if(reset2rx_client = '1' or eof_reset = '1') then
                    udp_pack_len_cntr_4 <= (others => '0');
                elsif(rx_client_clk_enbl = '1' and start_of_frame_array(initial_index + 52) = '1') then
          -- Load the counter with the UDP packet length and discount the #2-byte words till this point in time
          -- Counter Value = (UDP Pack Len/2) - 3. (#2-byte words already added to Checksum Calculation)
                    udp_pack_len_cntr_4_div2  := '0' & rxd_packed_16bits(15 downto 1);
                    udp_pack_len_cntr_4       <= udp_pack_len_cntr_4_div2-x"0003";   
                elsif(rx_client_clk_enbl = '1' and udp_pack_len_cntr_4 /= x"FFFF" and enable_udp_hdr_sum_4 = '1' and pack_high_1_pack_low_0 = '1') then
                    udp_pack_len_cntr_4 <= udp_pack_len_cntr_4-x"0001";
                end if;
            end if;
        end process;

        udp_len_is_odd_4  <= save_udp_hdr_length_4(0);
        udp_eof_reached_4 <= '1' when ((udp_pack_len_cntr_4 = x"0001" and udp_len_is_odd_4 = '0') or (udp_pack_len_cntr_4 = x"0000" and udp_len_is_odd_4 = '1')) 
                             else '0'; 

        ENABLE_UDP_HEADER_SUM_4_PROCESS: process (RX_CLIENT_CLK) -- yes vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_udp_hdr_sum_4  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 35) = '1') then
                            enable_udp_hdr_sum_4  <= '1';
                        elsif((udp_eof_reached_4 = '1' and pack_high_1_pack_low_0 = '1') or start_of_frame_d1 = '0') then
                            enable_udp_hdr_sum_4  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SAVE_TCP_LENGTH_1_PROCESS: process (RX_CLIENT_CLK) -- no vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    save_tcp_length_1  <= (others => '0');
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 18) = '1') then
                            save_tcp_length_1  <= std_logic_vector(rxd_packed_16bits - X"0014");
                        elsif(eof_reset = '1') then
                            save_tcp_length_1  <= (others => '0');
                        end if;
                    end if;
                end if;
            end if;
        end process;

        tcp_pack_len_cntr_1_process: process(rx_client_clk)
            variable tcp_pack_len_cntr_1_div2 : unsigned(15 downto 0);
        begin
            if(rising_edge(rx_client_clk)) then
                if(reset2rx_client = '1' or eof_reset = '1') then
                    tcp_pack_len_cntr_1 <= (others => '1');
                elsif(rx_client_clk_enbl = '1' and start_of_frame_array(initial_index + 18) = '1') then
                    tcp_pack_len_cntr_1_div2  := '0' & rxd_packed_16bits(15 downto 1);
                    tcp_pack_len_cntr_1       <= tcp_pack_len_cntr_1_div2-x"0004";   
                elsif(rx_client_clk_enbl = '1' and tcp_pack_len_cntr_1 /= x"FFFF" and enable_tcp_hdr_sum_1 = '1' and pack_high_1_pack_low_0 = '1') then
                    tcp_pack_len_cntr_1 <= tcp_pack_len_cntr_1-x"0001";
                end if;
            end if;
        end process;

        tcp_len_is_odd_1  <= save_tcp_length_1(0);
        tcp_eof_reached_1 <= '1' when ((tcp_pack_len_cntr_1 = x"0001" and tcp_len_is_odd_1 = '0') or (tcp_pack_len_cntr_1 = x"0000" and tcp_len_is_odd_1 = '1')) 
                             else '0'; 

        ENABLE_TCP_HEADER_SUM_1_PROCESS: process (RX_CLIENT_CLK) -- no vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_tcp_hdr_sum_1  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 23) = '1') then
                            enable_tcp_hdr_sum_1  <= '1';
                        elsif((tcp_eof_reached_1 = '1' and pack_high_1_pack_low_0 = '1') or start_of_frame_d1 = '0') then
                            enable_tcp_hdr_sum_1  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_TCP_HDR_1_PROCESS: process (RX_CLIENT_CLK) -- no vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    tcp_header_sum_1  <=(others => '0');
                    tcp_header_csum_1_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            tcp_header_csum_1_ok <= '0';
                        elsif ((tcp_header_sum_1(15 downto 0) + unsigned(save_tcp_length_1)) = X"FFFF" and tcp_header_sum_1(16) = '0' and enable_tcp_hdr_sum_1 = '0') then
                            tcp_header_csum_1_ok <= '1';
                        elsif ((tcp_header_sum_1(15 downto 0) + unsigned(save_tcp_length_1)) = X"FFFE" and tcp_header_sum_1(16) = '1' and enable_tcp_hdr_sum_1 = '0') then
                            tcp_header_csum_1_ok <= '1';
                        else
                            tcp_header_csum_1_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            tcp_header_sum_1  <=(others => '0');
                        elsif (enable_tcp_hdr_sum_1 = '1' and pack_high_1_pack_low_0 = '1') then
                            if (start_of_frame_array(initial_index + 24) = '1') then -- mask Time to live filed from protocol in Ip header
                                tcp_header_sum_1(16 downto 0)  <= ('0'&tcp_header_sum_1(15 downto 0)) + ("000000000"&rxd_packed_16bits(7 downto 0));
                            elsif (start_of_frame_array(initial_index + 26) = '1') then -- mask IP header csum
                                tcp_header_sum_1(16 downto 0)  <= ('0'&tcp_header_sum_1(15 downto 0)) + ("00000000000000000");
                            elsif(tcp_eof_reached_1 = '1' and tcp_len_is_odd_1 = '1') then
                                tcp_header_sum_1(16 downto 0)  <= ('0' & tcp_header_sum_1(15 downto 0)) + (rxd_packed_16bits(15 downto 8) & x"00");
                            else
                                tcp_header_sum_1(16 downto 0)  <= ('0'&tcp_header_sum_1(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                            end if;
                        elsif (enable_tcp_hdr_sum_1 = '1' and pack_high_1_pack_low_0 = '0') then
                            tcp_header_sum_1(16 downto 0)  <= ('0'&tcp_header_sum_1(15 downto 0)) + (X"0000"&tcp_header_sum_1(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SAVE_TCP_LENGTH_2_PROCESS: process (RX_CLIENT_CLK) -- yes vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    save_tcp_length_2  <= (others => '0');
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 22) = '1') then
                            save_tcp_length_2  <= std_logic_vector(rxd_packed_16bits - X"0014");
                        elsif(eof_reset = '1') then
                            save_tcp_length_2  <= (others => '0');
                        end if;
                    end if;
                end if;
            end if;
        end process;

        tcp_pack_len_cntr_2_process: process(rx_client_clk)
            variable tcp_pack_len_cntr_2_div2 : unsigned(15 downto 0);
        begin
            if(rising_edge(rx_client_clk)) then
                if(reset2rx_client = '1' or eof_reset = '1') then
                    tcp_pack_len_cntr_2 <= (others => '1');
                elsif(rx_client_clk_enbl = '1' and start_of_frame_array(initial_index + 22) = '1') then
                    tcp_pack_len_cntr_2_div2  := '0' & rxd_packed_16bits(15 downto 1);
                    tcp_pack_len_cntr_2       <= tcp_pack_len_cntr_2_div2-x"0004";   
                elsif(rx_client_clk_enbl = '1' and tcp_pack_len_cntr_2 /= x"FFFF" and enable_tcp_hdr_sum_2 = '1' and pack_high_1_pack_low_0 = '1') then
                    tcp_pack_len_cntr_2 <= tcp_pack_len_cntr_2-x"0001";
                end if;
            end if;
        end process;

        tcp_len_is_odd_2  <= save_tcp_length_2(0);
        tcp_eof_reached_2 <= '1' when ((tcp_pack_len_cntr_2 = x"0001" and tcp_len_is_odd_2 = '0') or (tcp_pack_len_cntr_2 = x"0000" and tcp_len_is_odd_2 = '1')) 
                             else '0'; 

        ENABLE_TCP_HEADER_SUM_2_PROCESS: process (RX_CLIENT_CLK) -- yes vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_tcp_hdr_sum_2  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 27) = '1') then
                            enable_tcp_hdr_sum_2  <= '1';
                        elsif((tcp_eof_reached_2 = '1' and pack_high_1_pack_low_0 = '1') or start_of_frame_d1 = '0') then
                            enable_tcp_hdr_sum_2  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_TCP_HDR_2_PROCESS: process (RX_CLIENT_CLK) -- yes vlan no snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    tcp_header_sum_2  <=(others => '0');
                    tcp_header_csum_2_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            tcp_header_csum_2_ok <= '0';
                        elsif ((tcp_header_sum_2(15 downto 0) + unsigned(save_tcp_length_2)) = X"FFFF" and tcp_header_sum_2(16) = '0' and enable_tcp_hdr_sum_2 = '0') then
                            tcp_header_csum_2_ok <= '1';
                        elsif ((tcp_header_sum_2(15 downto 0) + unsigned(save_tcp_length_2)) = X"FFFE" and tcp_header_sum_2(16) = '1' and enable_tcp_hdr_sum_2 = '0') then
                            tcp_header_csum_2_ok <= '1';
                        else
                            tcp_header_csum_2_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            tcp_header_sum_2  <=(others => '0');
                        elsif (enable_tcp_hdr_sum_2 = '1' and pack_high_1_pack_low_0 = '1') then
                            if (start_of_frame_array(initial_index + 28) = '1') then -- mask Time to live filed from protocol in Ip header
                                tcp_header_sum_2(16 downto 0)  <= ('0'&tcp_header_sum_2(15 downto 0)) + ("000000000"&rxd_packed_16bits(7 downto 0));
                            elsif (start_of_frame_array(initial_index + 30) = '1') then -- mask IP header csum
                                tcp_header_sum_2(16 downto 0)  <= ('0'&tcp_header_sum_2(15 downto 0)) + ("00000000000000000");
                            elsif(tcp_eof_reached_2 = '1' and tcp_len_is_odd_2 = '1') then
                                tcp_header_sum_2(16 downto 0)  <= ('0' & tcp_header_sum_2(15 downto 0)) + (rxd_packed_16bits(15 downto 8) & x"00");
                            else
                                tcp_header_sum_2(16 downto 0)  <= ('0'&tcp_header_sum_2(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                            end if;
                        elsif (enable_tcp_hdr_sum_2 = '1' and pack_high_1_pack_low_0 = '0') then
                            tcp_header_sum_2(16 downto 0)  <= ('0'&tcp_header_sum_2(15 downto 0)) + (X"0000"&tcp_header_sum_2(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SAVE_TCP_LENGTH_3_PROCESS: process (RX_CLIENT_CLK) -- no vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    save_tcp_length_3  <= (others => '0');
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 26) = '1') then
                            save_tcp_length_3  <= std_logic_vector(rxd_packed_16bits - X"0014");
                        elsif(eof_reset = '1') then
                            save_tcp_length_3  <= (others => '0');
                        end if;
                    end if;
                end if;
            end if;
        end process;

        tcp_pack_len_cntr_3_process: process(rx_client_clk)
            variable tcp_pack_len_cntr_3_div2 : unsigned(15 downto 0);
        begin
            if(rising_edge(rx_client_clk)) then
                if(reset2rx_client = '1' or eof_reset = '1') then
                    tcp_pack_len_cntr_3 <= (others => '1');
                elsif(rx_client_clk_enbl = '1' and start_of_frame_array(initial_index + 26) = '1') then
                    tcp_pack_len_cntr_3_div2  := '0' & rxd_packed_16bits(15 downto 1);
                    tcp_pack_len_cntr_3       <= tcp_pack_len_cntr_3_div2-x"0004";   
                elsif(rx_client_clk_enbl = '1' and tcp_pack_len_cntr_3 /= x"FFFF" and enable_tcp_hdr_sum_3 = '1' and pack_high_1_pack_low_0 = '1') then
                    tcp_pack_len_cntr_3 <= tcp_pack_len_cntr_3-x"0001";
                end if;
            end if;
        end process;

        tcp_len_is_odd_3  <= save_tcp_length_3(0);
        tcp_eof_reached_3 <= '1' when ((tcp_pack_len_cntr_3 = x"0001" and tcp_len_is_odd_3 = '0') or (tcp_pack_len_cntr_3 = x"0000" and tcp_len_is_odd_3 = '1')) 
                             else '0'; 

        ENABLE_TCP_HEADER_SUM_3_PROCESS: process (RX_CLIENT_CLK) -- no vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_tcp_hdr_sum_3  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 31) = '1') then
                            enable_tcp_hdr_sum_3  <= '1';
                        elsif((tcp_eof_reached_3 = '1' and pack_high_1_pack_low_0 = '1') or start_of_frame_d1 = '0') then
                            enable_tcp_hdr_sum_3  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_TCP_HDR_3_PROCESS: process (RX_CLIENT_CLK) -- no vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    tcp_header_sum_3  <=(others => '0');
                    tcp_header_csum_3_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            tcp_header_csum_3_ok <= '0';
                        elsif ((tcp_header_sum_3(15 downto 0) + unsigned(save_tcp_length_3)) = X"FFFF" and tcp_header_sum_3(16) = '0' and
                        enable_tcp_hdr_sum_3 = '0') then
                            tcp_header_csum_3_ok <= '1';
                        elsif ((tcp_header_sum_3(15 downto 0) + unsigned(save_tcp_length_3)) = X"FFFE" and tcp_header_sum_3(16) = '1' and
                        enable_tcp_hdr_sum_3 = '0') then
                            tcp_header_csum_3_ok <= '1';
                        else
                            tcp_header_csum_3_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            tcp_header_sum_3  <=(others => '0');
                        elsif (enable_tcp_hdr_sum_3 = '1' and pack_high_1_pack_low_0 = '1') then
                            if (start_of_frame_array(initial_index + 32) = '1') then -- mask Time to live filed from protocol in Ip header
                                tcp_header_sum_3(16 downto 0)  <= ('0'&tcp_header_sum_3(15 downto 0)) + ("000000000"&rxd_packed_16bits(7 downto 0));
                            elsif (start_of_frame_array(initial_index + 34) = '1') then -- mask IP header csum
                                tcp_header_sum_3(16 downto 0)  <= ('0'&tcp_header_sum_3(15 downto 0)) + ("00000000000000000");
                            elsif(tcp_eof_reached_3 = '1' and tcp_len_is_odd_3 = '1') then
                                tcp_header_sum_3(16 downto 0)  <= ('0' & tcp_header_sum_3(15 downto 0)) + (rxd_packed_16bits(15 downto 8) & x"00");
                            else
                                tcp_header_sum_3(16 downto 0)  <= ('0'&tcp_header_sum_3(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                            end if;
                        elsif (enable_tcp_hdr_sum_3 = '1' and pack_high_1_pack_low_0 = '0') then
                            tcp_header_sum_3(16 downto 0)  <= ('0'&tcp_header_sum_3(15 downto 0)) + (X"0000"&tcp_header_sum_3(16));

                        end if;
                    end if;
                end if;
            end if;
        end process;

        SAVE_TCP_LENGTH_4_PROCESS: process (RX_CLIENT_CLK) -- yes vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    save_tcp_length_4  <= (others => '0');
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 30) = '1') then
                            save_tcp_length_4  <= std_logic_vector(rxd_packed_16bits - X"0014");
                        elsif(eof_reset = '1') then
                            save_tcp_length_4  <= (others => '0');
                        end if;
                    end if;
                end if;
            end if;
        end process;

        tcp_pack_len_cntr_4_process: process(rx_client_clk)
            variable tcp_pack_len_cntr_4_div2 : unsigned(15 downto 0);
        begin
            if(rising_edge(rx_client_clk)) then
                if(reset2rx_client = '1' or eof_reset = '1') then
                    tcp_pack_len_cntr_4 <= (others => '1');
                elsif(rx_client_clk_enbl = '1' and start_of_frame_array(initial_index + 30) = '1') then
                    tcp_pack_len_cntr_4_div2  := '0' & rxd_packed_16bits(15 downto 1);
                    tcp_pack_len_cntr_4       <= tcp_pack_len_cntr_4_div2-x"0004";   
                elsif(rx_client_clk_enbl = '1' and tcp_pack_len_cntr_4 /= x"FFFF" and enable_tcp_hdr_sum_4 = '1' and pack_high_1_pack_low_0 = '1') then
                    tcp_pack_len_cntr_4 <= tcp_pack_len_cntr_4-x"0001";
                end if;
            end if;
        end process;

        tcp_len_is_odd_4  <= save_tcp_length_4(0);
        tcp_eof_reached_4 <= '1' when ((tcp_pack_len_cntr_4 = x"0001" and tcp_len_is_odd_4 = '0') or (tcp_pack_len_cntr_4 = x"0000" and tcp_len_is_odd_4 = '1')) 
                             else '0'; 

        ENABLE_TCP_HEADER_SUM_4_PROCESS: process (RX_CLIENT_CLK) -- yes vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    enable_tcp_hdr_sum_4  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(initial_index + 35) = '1') then
                            enable_tcp_hdr_sum_4  <= '1';
                        elsif((tcp_eof_reached_4 = '1' and pack_high_1_pack_low_0 = '1') or start_of_frame_d1 = '0') then
                            enable_tcp_hdr_sum_4  <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        SUM_TCP_HDR_4_PROCESS: process (RX_CLIENT_CLK) -- yes vlan yes snap
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    tcp_header_sum_4  <=(others => '0');
                    tcp_header_csum_4_ok <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (eof_reset = '1') then
                            tcp_header_csum_4_ok <= '0';
                        elsif ((tcp_header_sum_4(15 downto 0) + unsigned(save_tcp_length_4)) = X"FFFF" and tcp_header_sum_4(16) = '0' and
                        enable_tcp_hdr_sum_4 = '0') then
                            tcp_header_csum_4_ok <= '1';
                        elsif ((tcp_header_sum_4(15 downto 0) + unsigned(save_tcp_length_4)) = X"FFFE" and tcp_header_sum_4(16) = '1' and
                        enable_tcp_hdr_sum_4 = '0') then
                            tcp_header_csum_4_ok <= '1';
                        else
                            tcp_header_csum_4_ok <= '0';
                        end if;

                        if (eof_reset = '1') then
                            tcp_header_sum_4  <=(others => '0');
                        elsif (enable_tcp_hdr_sum_4 = '1' and pack_high_1_pack_low_0 = '1') then
                            if (start_of_frame_array(initial_index + 36) = '1') then -- mask Time to live filed from protocol in Ip header
                                tcp_header_sum_4(16 downto 0)  <= ('0'&tcp_header_sum_4(15 downto 0)) + ("000000000"&rxd_packed_16bits(7 downto 0));
                            elsif (start_of_frame_array(initial_index + 38) = '1') then -- mask IP header csum
                                tcp_header_sum_4(16 downto 0)  <= ('0'&tcp_header_sum_4(15 downto 0)) + ("00000000000000000");
                            elsif(tcp_eof_reached_4 = '1' and tcp_len_is_odd_4 = '1') then
                                tcp_header_sum_4(16 downto 0)  <= ('0' & tcp_header_sum_4(15 downto 0)) + (rxd_packed_16bits(15 downto 8) & x"00");
                            else
                                tcp_header_sum_4(16 downto 0)  <= ('0'&tcp_header_sum_4(15 downto 0)) + ('0'&rxd_packed_16bits(15 downto 0));
                            end if;
                        elsif (enable_tcp_hdr_sum_4 = '1' and pack_high_1_pack_low_0 = '0') then
                            tcp_header_sum_4(16 downto 0)  <= ('0'&tcp_header_sum_4(15 downto 0)) + (X"0000"&tcp_header_sum_4(16));
                        end if;
                    end if;
                end if;
            end if;
        end process;

        CONTROL_16BIT_PACK_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    pack_high_1_pack_low_0  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (start_of_frame_array(1) = '1') then
                            pack_high_1_pack_low_0  <= '1';
                        else
                            pack_high_1_pack_low_0  <= not(pack_high_1_pack_low_0);
                        end if;
                    end if;
                end if;
            end if;
        end process;

        RXD_16BIT_PACK_PROCESS: process (RX_CLIENT_CLK)
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    rxd_packed_16bits  <= (others => '0');
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (pack_high_1_pack_low_0 = '1' and EMAC_CLIENT_RXD_VLD_LEGACY = '1') then
                            rxd_packed_16bits(15 downto 8) <= unsigned(EMAC_CLIENT_RXD_LEGACY);
                            rxd_packed_16bits(7 downto 0)  <= (others => '0');
                        elsif (pack_high_1_pack_low_0 = '0' and EMAC_CLIENT_RXD_VLD_LEGACY = '1') then
                            rxd_packed_16bits(7 downto 0)  <= unsigned(EMAC_CLIENT_RXD_LEGACY);
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -------------------------------------------------------------------------
    -- detect if the frame is a IPv4 Ethernet II frame with type 0800
    -------------------------------------------------------------------------

        DETECT_TYPE_0800 : process(RX_CLIENT_CLK)
    -- delay this check by one pipeline stage so we can detect vlan first valid by byte 22 when vlan
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_has_type_0800_d22   <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (frame_is_vlan_8100_d15 = '0') then -- no vlan
                            if (((rx_data_words_array(1)(7 downto 0) & rx_data_words_array(1)(15 downto 8)) = X"0800") and start_of_frame_array(initial_index + 17) = '1') then
                                frame_has_type_0800_d22 <= '1';
                            elsif (eof_reset = '1') then
                                frame_has_type_0800_d22 <= '0';
                            end if;
                        else -- vlan
                            if (((rx_data_words_array(1)(7 downto 0) & rx_data_words_array(1)(15 downto 8)) = X"0800") and start_of_frame_array(initial_index + 21) = '1') then
                                frame_has_type_0800_d22 <= '1';
                            elsif (eof_reset = '1') then
                                frame_has_type_0800_d22 <= '0';
                            end if;
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -------------------------------------------------------------------------
    -- detect if the frame has a valid length field
    -------------------------------------------------------------------------

        DETECT_VALID_LENGTH_FIELD : process(RX_CLIENT_CLK)
    -- delay this check by one pipeline stage so we can detect vlan first valid by byte 22 when vlan
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_has_valid_length_field_d22   <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (frame_is_vlan_8100_d15 = '0') then -- no vlan
                            if (((rx_data_words_array(1)(7 downto 0) & rx_data_words_array(1)(15 downto 8)) < X"0601") and
                            start_of_frame_array(initial_index + 17) = '1') then
                                frame_has_valid_length_field_d22 <= '1';
                            elsif (eof_reset = '1') then
                                frame_has_valid_length_field_d22 <= '0';
                            end if;
                        else -- vlan
                            if (((rx_data_words_array(1)(7 downto 0) & rx_data_words_array(1)(15 downto 8)) < X"0601") and
                            start_of_frame_array(initial_index + 21) = '1') then
                                frame_has_valid_length_field_d22 <= '1';
                            elsif (eof_reset = '1') then
                                frame_has_valid_length_field_d22 <= '0';
                            end if;
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -------------------------------------------------------------------------
    -- detect if the frame has an IPv4 protocol field value of 4
    -------------------------------------------------------------------------

        DETECT_IP_PROTO_FIELD : process(RX_CLIENT_CLK)
    -- delay this check by pipeline stages so we can detect snap first. valid by byte 31
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_is_ip_protocol_d31   <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (frame_is_vlan_8100_d15 = '0' and frame_is_snap_d30 = '0' and start_of_frame_array(initial_index + 30) = '1') then
              -- no vlan and no snap
                            if (((rx_data_words_array(4)(23 downto 20)) = X"4")) then
                                frame_is_ip_protocol_d31 <= '1';
                            end if;
                        elsif (frame_is_vlan_8100_d15 = '1' and frame_is_snap_d30 = '0' and start_of_frame_array(initial_index + 30) = '1') then
              -- yes vlan and no snap
                            if (((rx_data_words_array(3)(23 downto 20)) = X"4")) then
                                frame_is_ip_protocol_d31 <= '1';
                            end if;
                        elsif (frame_is_vlan_8100_d15 = '1' and frame_is_snap_d30 = '1' and start_of_frame_array(initial_index + 30) = '1') then
              -- yes vlan and yes snap
                            if (((rx_data_words_array(1)(23 downto 20)) = X"4")) then
                                frame_is_ip_protocol_d31 <= '1';
                            end if;
                        elsif (frame_is_vlan_8100_d15 = '0' and frame_is_snap_d30 = '1' and start_of_frame_array(initial_index + 30) = '1') then
              -- no vlan and yes snap
                            if (((rx_data_words_array(2)(23 downto 20)) = X"4")) then
                                frame_is_ip_protocol_d31 <= '1';
                            end if;
                        else
                            if (eof_reset = '1') then
                                frame_is_ip_protocol_d31 <= '0';
                            end if;
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -------------------------------------------------------------------------
    -- detect if the frame has an IPv4 header length field value of 5
    -------------------------------------------------------------------------

        DETECT_IP_HDR_LEN_FIELD : process(RX_CLIENT_CLK)
    -- delay this check by pipeline stages so we can detect snap first. valid by byte 31
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_has_ip_hdr_length_d31   <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (frame_is_vlan_8100_d15 = '0' and frame_is_snap_d30 = '0' and start_of_frame_array(initial_index + 30) = '1') then
              -- no vlan and no snap
                            if (((rx_data_words_array(4)(19 downto 16)) = X"5")) then
                                frame_has_ip_hdr_length_d31 <= '1';
                            end if;
                        elsif (frame_is_vlan_8100_d15 = '1' and frame_is_snap_d30 = '0' and start_of_frame_array(initial_index + 30) = '1') then
              -- yes vlan and no snap
                            if (((rx_data_words_array(3)(19 downto 16)) = X"5")) then
                                frame_has_ip_hdr_length_d31 <= '1';
                            end if;
                        elsif (frame_is_vlan_8100_d15 = '1' and frame_is_snap_d30 = '1' and start_of_frame_array(initial_index + 30) = '1') then
              -- yes vlan and yes snap
                            if (((rx_data_words_array(1)(19 downto 16)) = X"5")) then
                                frame_has_ip_hdr_length_d31 <= '1';
                            end if;
                        elsif (frame_is_vlan_8100_d15 = '0' and frame_is_snap_d30 = '1' and start_of_frame_array(initial_index + 30) = '1') then
              -- no vlan and yes snap
                            if (((rx_data_words_array(2)(19 downto 16)) = X"5")) then
                                frame_has_ip_hdr_length_d31 <= '1';
                            end if;
                        else
                            if (eof_reset = '1') then
                                frame_has_ip_hdr_length_d31 <= '0';
                            end if;
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -------------------------------------------------------------------------
    -- detect if the frame has a IPv4 fragments
    -------------------------------------------------------------------------

        DETECT_IP_FRAGS : process(RX_CLIENT_CLK)
    -- delay this check by pipeline stages so we can detect IP protocol and IP header length first. valid by byte 38
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_has_no_ip_frags_d38   <= '0';
                    frame_has_udp_protocol_d38  <= '0';
                    frame_has_tcp_protocol_d38  <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (frame_is_vlan_8100_d15 = '0' and frame_is_snap_d30 = '0' and frame_has_ip_hdr_length_d31= '1' and
                        frame_is_ip_protocol_d31 = '1' and start_of_frame_array(initial_index + 32) = '1') then -- no vlan and no snap
                            if (((rx_data_words_array(2)(5 downto 0)) = "000000") and ((rx_data_words_array(2)(15 downto 7)) = "000000000")) then
                -- skip bit 6 which is don't framement flag which is allowed to be set
                                frame_has_no_ip_frags_d38 <= '1';
                            end if;
                            if (((rx_data_words_array(2)(31 downto 24)) = X"11")) then
                                frame_has_udp_protocol_d38 <= '1';
                                frame_has_tcp_protocol_d38 <= '0';
                            end if;
                            if (((rx_data_words_array(2)(31 downto 24)) = X"06")) then
                                frame_has_udp_protocol_d38 <= '0';
                                frame_has_tcp_protocol_d38 <= '1';
                            end if;
                        elsif (frame_is_vlan_8100_d15 = '1' and frame_is_snap_d30 = '0' and frame_has_ip_hdr_length_d31= '1' and
                        frame_is_ip_protocol_d31 = '1' and start_of_frame_array(initial_index + 32) = '1') then -- yes vlan and no snap
                            if (((rx_data_words_array(1)(5 downto 0)) = "000000") and ((rx_data_words_array(1)(15 downto 7)) = "000000000")) then
                -- skip bit 6 which is don't framement flag which is allowed to be set
                                frame_has_no_ip_frags_d38 <= '1';
                            end if;
                            if (((rx_data_words_array(1)(31 downto 24)) = X"11")) then
                                frame_has_udp_protocol_d38 <= '1';
                                frame_has_tcp_protocol_d38 <= '0';
                            end if;
                            if (((rx_data_words_array(1)(31 downto 24)) = X"06")) then
                                frame_has_udp_protocol_d38 <= '0';
                                frame_has_tcp_protocol_d38 <= '1';
                            end if;
                        elsif (frame_is_vlan_8100_d15 = '1' and frame_is_snap_d30 = '1' and frame_has_ip_hdr_length_d31= '1' and
                        frame_is_ip_protocol_d31 = '1' and start_of_frame_array(initial_index + 40) = '1') then -- yes vlan and yes snap
                            if (((rx_data_words_array(1)(5 downto 0)) = "000000") and ((rx_data_words_array(1)(15 downto 7)) = "000000000")) then
                -- skip bit 6 which is don't framement flag which is allowed to be set
                                frame_has_no_ip_frags_d38 <= '1';
                            end if;
                            if (((rx_data_words_array(1)(31 downto 24)) = X"11")) then
                                frame_has_udp_protocol_d38 <= '1';
                                frame_has_tcp_protocol_d38 <= '0';
                            end if;
                            if (((rx_data_words_array(1)(31 downto 24)) = X"06")) then
                                frame_has_udp_protocol_d38 <= '0';
                                frame_has_tcp_protocol_d38 <= '1';
                            end if;
                        elsif (frame_is_vlan_8100_d15 = '0' and frame_is_snap_d30 = '1' and frame_has_ip_hdr_length_d31= '1' and
                        frame_is_ip_protocol_d31 = '1' and start_of_frame_array(initial_index + 36) = '1') then -- no vlan and yes snap
                            if (((rx_data_words_array(1)(5 downto 0)) = "000000") and ((rx_data_words_array(1)(15 downto 7)) = "000000000")) then
                -- skip bit 6 which is don't framement flag which is allowed to be set
                                frame_has_no_ip_frags_d38 <= '1';
                            end if;
                            if (((rx_data_words_array(1)(31 downto 24)) = X"11")) then
                                frame_has_udp_protocol_d38 <= '1';
                                frame_has_tcp_protocol_d38 <= '0';
                            end if;
                            if (((rx_data_words_array(1)(31 downto 24)) = X"06")) then
                                frame_has_udp_protocol_d38 <= '0';
                                frame_has_tcp_protocol_d38 <= '1';
                            end if;
                        else
                            if (eof_reset = '1') then
                                frame_has_no_ip_frags_d38 <= '0';
                                frame_has_udp_protocol_d38 <= '0';
                                frame_has_tcp_protocol_d38 <= '0';
                            end if;
                        end if;
                    end if;
                end if;
            end if;
        end process;

    -------------------------------------------------------------------------
    -- detect if the frame has a IPv4 Ethernet SNAP frame with type 0800
    -------------------------------------------------------------------------

        DETECT_SNAP : process(RX_CLIENT_CLK)
    -- delay this check by one pipeline stage so we can detect vlan first valid by byte 30 when vlan
        begin
            if rising_edge(RX_CLIENT_CLK) then
                if RESET2RX_CLIENT = '1' then
                    frame_is_snap_d30   <= '0';
                else
                    if (RX_CLIENT_CLK_ENBL = '1') then
                        if (frame_is_vlan_8100_d15 = '0') then -- no vlan
                            if ((rx_data_words_array(3)(31 downto 16) = X"AAAA") and
                            (rx_data_words_array(2)(31 downto 0) =  X"00000003") and
                            (rx_data_words_array(1)(15 downto 0) =  X"0008") and
                            start_of_frame_array(initial_index + 25) = '1') and (frame_has_valid_length_field_d22 = '1') then
                                frame_is_snap_d30 <= '1';
                            elsif (eof_reset = '1') then
                                frame_is_snap_d30 <= '0';
                            end if;
                        else -- vlan
                            if ((rx_data_words_array(3)(31 downto 16) = X"AAAA") and
                            (rx_data_words_array(2)(31 downto 0) =  X"00000003") and
                            (rx_data_words_array(1)(15 downto 0) =  X"0008") and
                            start_of_frame_array(initial_index + 29) = '1') and (frame_has_valid_length_field_d22 = '1') then
                                frame_is_snap_d30 <= '1';
                            elsif (eof_reset = '1') then
                                frame_is_snap_d30 <= '0';
                            end if;
                        end if;
                    end if;
                end if;
            end if;
        end process;
    end generate YES_FULL_CSUM_OFFLOAD;

  -------------------------------------------------------------------------
  -- Synchronize gray encoded last processed pointer from AXIStream clock
  -- domain to the receive client clock domain.
  -------------------------------------------------------------------------
    SYNC_RXS_LAST_READ_GRAY_PROCESS: for i in 35 downto 0 generate
        SYNC_RXS_LAST_READ_GRAY: sync_block
        port map (
                     clk       => RX_CLIENT_CLK,
                     reset     => RESET2RX_CLIENT,
                     data_in   => AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY(i),
                     data_out  => sync_rxs_mem_last_read_out_ptr_gray_sync(i)
                 );
    end generate;

  -------------------------------------------------------------------------
  -- Convert gray encoded last processed pointer back to binary encoded
  -------------------------------------------------------------------------
    rxclclk_rxs_mem_last_read_out_ptr <= unsigned(gray_to_bin(sync_rxs_mem_last_read_out_ptr_gray_sync));

  -------------------------------------------------------------------------
  -- Register binary encoded last processed pointer from local link
  -- interface
  -------------------------------------------------------------------------
    RX_CL_CLK_REG_RXS_LAST_READ_PROCESS: process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                rxclclk_rxs_mem_last_read_out_ptr_d1  <= (others => '0');
            else
                rxclclk_rxs_mem_last_read_out_ptr_d1  <= rxclclk_rxs_mem_last_read_out_ptr;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- Synchronize gray encoded last processed pointer from AXIStream clock
  -- domain to the receive client clock domain.
  -------------------------------------------------------------------------
    SYNC_RXD_LAST_READ_GRAY_PROCESS: for i in 35 downto 0 generate
        SYNC_RXD_LAST_READ_GRAY: sync_block
        port map (
                     clk       => RX_CLIENT_CLK,
                     reset     => RESET2RX_CLIENT,
                     data_in   => AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY(i),
                     data_out  => sync_rxd_mem_last_read_out_ptr_gray_sync(i)
                 );
    end generate;

  -------------------------------------------------------------------------
  -- Convert gray encoded last processed pointer back to binary encoded
  -------------------------------------------------------------------------
    rxclclk_rxd_mem_last_read_out_ptr <= gray_to_bin(sync_rxd_mem_last_read_out_ptr_gray_sync);

  -------------------------------------------------------------------------
  -- Register binary encoded last processed pointer from local link
  -- interface
  -------------------------------------------------------------------------
    RX_CL_CLK_REG_RXD_LAST_READ_PROCESS: process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                rxclclk_rxd_mem_last_read_out_ptr_d1  <= (others => '0');
            else
                rxclclk_rxd_mem_last_read_out_ptr_d1  <= rxclclk_rxd_mem_last_read_out_ptr;
            end if;
        end if;
    end process;

  -----------------------------------------------------------------------------

    rxs_status_word_2               <= X"00000" & multicast_addr_upper_d10;
    rxs_status_word_3               <= X"0" & multicast_addr_lower_d10;
    rxs_status_word_4               <= X"0" & statistics_vector & receive_checksum_status & frame_is_broadcast_d10 &
                                       frame_is_ip_multicast_d4 & frame_is_multicast_d10;
    rxs_status_word_5               <= X"0" & bytes_12_and_13_d19 & raw_checksum;
    rxs_status_word_6_cmb(35 downto 16) <= X"0" & bytes_14_and_15_d19;

    RX_CL_CLK_VLAN_ADDR         <= (others => '0');
    RX_CL_CLK_VLAN_BRAM_EN_A    <= '0';

  -------------------------------------------------------------------------
  -- Generate variable width address masks for checking memory pointers
  -------------------------------------------------------------------------
    RXD_GEN_MASK: for I in C_RXD_MEM_ADDR_WIDTH downto 0 generate
        rxd_mem_full_mask(I) <= '1';
        rxd_mem_empty_mask(I)  <= '0';
    end generate;

    rxd_mem_one_mask            <= unsigned(rxd_mem_empty_mask) + 1;
    rxd_mem_two_mask            <= unsigned(rxd_mem_empty_mask) + 2;
    rxd_mem_full_mask_minus_one <= rxd_mem_full_mask - 1;

    RXS_GEN_MASK: for I in C_RXS_MEM_ADDR_WIDTH downto 0 generate
        rxs_mem_full_mask(I) <= '1';
        rxs_mem_empty_mask(I)  <= '0';
    end generate;

    rxs_mem_one_mask            <= rxs_mem_empty_mask + 1;
    rxs_mem_two_mask            <= rxs_mem_empty_mask + 2;
    rxs_mem_three_mask          <= rxs_mem_empty_mask + 3;
    rxs_mem_four_mask           <= rxs_mem_empty_mask + 4;
    rxs_mem_full_mask_minus_one <= rxs_mem_full_mask - 1;

    zero_extend_rxd_mask36      <= (others => '0');
    zero_extend_rxs_mask36      <= (others => '0');

  -------------------------------------------------------------------------
  -- pack the 8 bit wide client receive data into 32 bit wide
  -------------------------------------------------------------------------

    RX_DATA_8_TO_32_PACK : process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                rx_data_packed_word      <= (others => '0');
                rx_data_vld_packed_word  <= (others => '0');
                rx_data_packed_state     <= (others => '0');
                rx_data_packed_ready     <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (EMAC_CLIENT_RXD_VLD_LEGACY = '1') then -- word full and ready to use
                        if (rx_data_packed_state = "11") then
                            rx_data_packed_state <= (others => '0');
                            rx_data_packed_ready <= '1';
                        else
                            rx_data_packed_state <= std_logic_vector(unsigned(rx_data_packed_state) + 1);
                            rx_data_packed_ready <= '0';
                        end if;
                        if (rx_data_packed_state = "00") then
                            rx_data_vld_packed_word(3)        <= EMAC_CLIENT_RXD_VLD_LEGACY;
                            rx_data_packed_word(31 downto 24) <= EMAC_CLIENT_RXD_LEGACY;
                        elsif(rx_data_packed_state = "01") then
                            rx_data_vld_packed_word(3 downto 2) <= EMAC_CLIENT_RXD_VLD_LEGACY & rx_data_vld_packed_word(3);
                            rx_data_packed_word(31 downto 16)   <= EMAC_CLIENT_RXD_LEGACY & rx_data_packed_word(31 downto 24);
                        elsif(rx_data_packed_state = "10") then
                            rx_data_vld_packed_word(3 downto 1) <= EMAC_CLIENT_RXD_VLD_LEGACY & rx_data_vld_packed_word(3 downto 2);
                            rx_data_packed_word(31 downto 8)    <= EMAC_CLIENT_RXD_LEGACY     & rx_data_packed_word(31 downto 16);
                        elsif(rx_data_packed_state = "11") then
                            rx_data_vld_packed_word(3 downto 0) <= EMAC_CLIENT_RXD_VLD_LEGACY & rx_data_vld_packed_word(3 downto 1);
                            rx_data_packed_word(31 downto 0)    <= EMAC_CLIENT_RXD_LEGACY     & rx_data_packed_word(31 downto 8);
                        end if;
                    elsif (EMAC_CLIENT_RXD_VLD_LEGACY = '0' and rx_data_valid_array(1)(0) = '1') then
                        if(rx_data_packed_state = "01") then
                            rx_data_vld_packed_word(3 downto 0) <= "000" & rx_data_vld_packed_word(3);
                            rx_data_packed_word(31 downto 0)    <= "000000000000000000000000" & rx_data_packed_word(31 downto 24);
                            rx_data_packed_ready <= '1';
                            rx_data_packed_state     <= (others => '0');
                        elsif(rx_data_packed_state = "10") then
                            rx_data_vld_packed_word(3 downto 0) <= "00" & rx_data_vld_packed_word(3 downto 2);
                            rx_data_packed_word(31 downto 0)    <= "0000000000000000" & rx_data_packed_word(31 downto 16);
                            rx_data_packed_ready <= '1';
                            rx_data_packed_state     <= (others => '0');
                        elsif(rx_data_packed_state = "11") then
                            rx_data_vld_packed_word(3 downto 0) <= '0' & rx_data_vld_packed_word(3 downto 1);
                            rx_data_packed_word(31 downto 0)    <= "00000000" & rx_data_packed_word(31 downto 8);
                            rx_data_packed_ready <= '1';
                            rx_data_packed_state     <= (others => '0');
                        else
                            rx_data_packed_word      <= (others => '0');
                            rx_data_vld_packed_word  <= (others => '0');
                            rx_data_packed_state     <= (others => '0');
                            rx_data_packed_ready     <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- calculate the partial checksum or not
  -------------------------------------------------------------------------

    INCLUDE_RX_CSUM: if(C_RXCSUM = 1) generate
        signal emacClientRxdLegacy_d1    : std_logic_vector(7 downto 0);
        signal rxd16bits                 : std_logic_vector(15 downto 0);
        signal emacClientRxdVldLegacy_d1 : std_logic;
        signal emacClientRxdVldWord      : std_logic;
    begin
        process(RX_CLIENT_CLK)
        begin
            if(rising_edge(RX_CLIENT_CLK)) then
                if(RESET2RX_CLIENT='1') then
                    emacClientRxdLegacy_d1   <= (others => '0');
                    emacClientRxdVldWord<= '0';
                else
                    if(RX_CLIENT_CLK_ENBL='1') then
                        emacClientRxdLegacy_d1   <= EMAC_CLIENT_RXD_LEGACY;
                        emacClientRxdVldLegacy_d1<= EMAC_CLIENT_RXD_VLD_LEGACY;
                        if (EMAC_CLIENT_RXD_VLD_LEGACY = '1' or emacClientRxdVldLegacy_d1 = '1') then
                            emacClientRxdVldWord <= NOT(emacClientRxdVldWord);
                        else
                            emacClientRxdVldWord<= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        rxd16bits <= emacClientRxdLegacy_d1 & EMAC_CLIENT_RXD_LEGACY when EMAC_CLIENT_RXD_VLD_LEGACY = '1' else
                     emacClientRxdLegacy_d1 & X"00";

        I_RX_CSUM : rx_csum_if
        port map(
                    CLK       => RX_CLIENT_CLK,
                    CLK_ENBL  => RX_CLIENT_CLK_ENBL,
                    RST       => RESET2RX_CLIENT,
                    INTRFRMRST=> eof_reset,
                    CALC_ENBL => emacClientRxdVldLegacy_d1,
                    WORD_ENBL => emacClientRxdVldWord,
                    DATA_IN   => rxd16bits,
                    CSUM_VLD  => rxCsumVld,
                    CSUM      => rxCsum
                );
    end generate INCLUDE_RX_CSUM;

    EXCLUDE_RX_CSUM: if (not (C_RXCSUM = 1)) generate
    begin
        rxCsum <= (others => '0');
        rxCsumVld <= '0';
    end generate EXCLUDE_RX_CSUM;

  -------------------------------------------------------------------------
  -- save partial csum value once calculated
  -------------------------------------------------------------------------

    SAVE_PARTIAL_CSUM_VAL : process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                raw_checksum <= (others => '0');
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (eof_reset = '1') then -- clear at end of frame
                        raw_checksum <= (others => '0');
                    elsif (rxCsumVld = '1') then
                        raw_checksum <= rxCsum;
                    end if;
                end if;
            end if;
        end if;
    end process;

    -------------------------------------------------------------------------
    -- capture the statistics which is different for soft and hard TEMAC
    -------------------------------------------------------------------------

    frame_drop <= (EMAC_CLIENT_RX_STATS_VLD and not (SOFT_EMAC_CLIENT_RX_STATS(27)));

    CAPTURE_STATS : process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                statistics_vector <= (others => '0');
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (EMAC_CLIENT_RX_STATS_VLD = '1') then
                        statistics_vector(25 downto 22) <= SOFT_EMAC_CLIENT_RX_STATS(26 downto 23);
                        statistics_vector(21 downto 0) <= SOFT_EMAC_CLIENT_RX_STATS(21 downto 0);
                    end if;
                end if;
            end if;
        end if;

    end process;

  -------------------------------------------------------------------------
  -- count the number of bytes in the frame being received for 8 bit interface
  -------------------------------------------------------------------------

    COUNT_FRAME_RX_BYTES : process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                frame_length_bytes     <= (others => '0');
                frame_length_bytes_lat <= (others => '0');
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (end_of_frame_array(1) = '1') then -- clear at end of frame
                        frame_length_bytes <= (others => '0');
                    elsif (EMAC_CLIENT_RXD_VLD_LEGACY = '1') then
                        frame_length_bytes <= frame_length_bytes + 1;
                    end if;

                    if (end_of_frame_array(1) = '1') then
                        frame_length_bytes_lat <= frame_length_bytes;
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- save the good frame pulse so we can check it later
  -------------------------------------------------------------------------

    SAVE_GOOD_FRAME : process(RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                save_rx_goodframe   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (EMAC_CLIENT_RX_GOODFRAME_LEGACY = '1') then
                        save_rx_goodframe <= '1';
                    elsif (eof_reset = '1') then
                        save_rx_goodframe <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- save the bad frame pulse so we can check it later
  -------------------------------------------------------------------------

    SAVE_BAD_FRAME : process(RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                save_rx_badframe   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (EMAC_CLIENT_RX_BADFRAME_LEGACY = '1') then
                        save_rx_badframe <= '1';
                    elsif (eof_reset = '1') then
                        save_rx_badframe <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- check for not enough rxs memory
  -------------------------------------------------------------------------

    CHECK_RXS_MEM_AVAIL : process(RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                not_enough_rxs_memory   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
          -- rxs_mem_last_read_out_ptr_cmb being read out of rxs memory during state END_OF_FRAME_CHECK_GOOD_BAD
                    if (rxs_mem_addr_cntr   = rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0) or
                    rxs_mem_addr_cntr+1 = rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0) or
                    rxs_mem_addr_cntr+2 = rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0) or
                    rxs_mem_addr_cntr+3 = rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0) or
                    rxs_mem_addr_cntr+4 = rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0) or
                    rxs_mem_addr_cntr+5 = rxclclk_rxs_mem_last_read_out_ptr_d1(C_RXS_MEM_ADDR_WIDTH downto 0)) then
                        not_enough_rxs_memory <= '1';
                    else
                        not_enough_rxs_memory <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- create a pipeline of receive data, receive data valid, start of frame
  -- end of frame
  -------------------------------------------------------------------------

    PIPE_RX_INPUTS_4 : process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                rx_data_words_array   <= (others => (others => '0'));
                rx_data_valid_array   <= (others => (others => '0'));
                end_of_frame_array    <= (others => '0');
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    end_of_frame_array (1)      <= start_of_frame_d1 and not(EMAC_CLIENT_RXD_VLD_LEGACY);
                    if (rx_data_packed_ready = '1') then
                        rx_data_words_array (1)     <= rx_data_packed_word;
                        rx_data_valid_array (1)     <= rx_data_vld_packed_word;
                    end if;
                    for i in 1 to 3 loop
                        end_of_frame_array (i+1)     <= end_of_frame_array (i);
                        if (rx_data_packed_ready = '1') then
                            rx_data_words_array (i+1)  <= rx_data_words_array (i);
                            rx_data_valid_array (i+1)  <= rx_data_valid_array (i);
                        end if;
                    end loop;
                end if;
            end if;
        end if;
    end process;

    PIPE_RX_INPUTS_100_12 : process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                start_of_frame_d1     <= '0';
                start_of_frame_array  <= (others => '0');
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    start_of_frame_d1           <= EMAC_CLIENT_RXD_VLD_LEGACY;
                    start_of_frame_array (1)    <= EMAC_CLIENT_RXD_VLD_LEGACY and not(start_of_frame_d1);
                    for i in 1 to 51 loop
                        start_of_frame_array (i+1)   <= start_of_frame_array (i);
                    end loop;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the destination address is broadcast
  -------------------------------------------------------------------------

    DETECT_BROADCAST : process(RX_CLIENT_CLK) -- valid by byte 10
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                frame_is_broadcast_d10   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (rx_data_words_array(1)(15 downto 0)  = X"FFFF" and
                    rx_data_words_array(2)(31 downto 0) = X"FFFFFFFF" and
                    start_of_frame_array(initial_index + 9) = '1') then
                        frame_is_broadcast_d10 <= '1';
                    elsif (eof_reset = '1') then
                        frame_is_broadcast_d10 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the destination address is IP multicast
  -------------------------------------------------------------------------

    DETECT_IP_MULTICAST : process(RX_CLIENT_CLK) -- valid by byte 4
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                frame_is_ip_multicast_d4   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (rx_data_packed_word(31 downto 24) = X"5E" and
                    rx_data_packed_word(23 downto 16) = X"00" and
                    rx_data_packed_word(15 downto 8)  = X"01" and
                    start_of_frame_array(initial_index + 3) = '1') then
                        frame_is_ip_multicast_d4 <= '1';
                    elsif (eof_reset = '1') then
                        frame_is_ip_multicast_d4 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the destination address is any multicast
  -------------------------------------------------------------------------

    DETECT_MULTICAST : process(RX_CLIENT_CLK) -- valid by byte 10
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                frame_is_multicast_d10   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (rx_data_words_array(2)(0) = '1' and
                    not((rx_data_words_array(1)(15 downto 0)  = X"FFFF")and
                    (rx_data_words_array(2)(31 downto 0) = X"FFFFFFFF"))and
                    start_of_frame_array(initial_index + 9) = '1') then
                        frame_is_multicast_d10 <= '1';
                    elsif (eof_reset = '1') then
                        frame_is_multicast_d10 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- save the destination (multicast) address for AXIStream status words
  -------------------------------------------------------------------------

    SAVE_DEST_ADDR : process(RX_CLIENT_CLK) -- valid by byte 10
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                multicast_addr_upper_d10   <= (others => '0');
                multicast_addr_lower_d10   <= (others => '0');
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (start_of_frame_array(initial_index + 9) = '1') then
                        multicast_addr_upper_d10 <= rx_data_words_array(1)(15 downto 0);
                        multicast_addr_lower_d10 <= rx_data_words_array(2)(31 downto 0);
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- save the bytes 12 thru 15 for AXIStream status words
  -------------------------------------------------------------------------

    SAVE_BYTES_12_TO_14 : process(RX_CLIENT_CLK) -- valid by byte 19
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                bytes_12_and_13_d19   <= (others => '0');
                bytes_14_and_15_d19   <= (others => '0');
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (start_of_frame_array(initial_index + 18) = '1') then
                        bytes_12_and_13_d19 <= rx_data_words_array(1)(15 downto 0);
                        bytes_14_and_15_d19 <= rx_data_words_array(1)(31 downto 16);
                    end if;
                end if;
            end if;
        end if;
    end process;

    -------------------------------------------------------------------------
    -- detect if the frame is a VLAN with type 8100
    -------------------------------------------------------------------------

    DETECT_VLAN_8100 : process(RX_CLIENT_CLK) -- valid by byte 15
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                frame_is_vlan_8100_d15   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = X"8100") and start_of_frame_array(initial_index + 14) = '1') then
                        frame_is_vlan_8100_d15 <= '1';
                    elsif (eof_reset = '1') then
                        frame_is_vlan_8100_d15 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a first VLAN tag with type TPID 0
  -------------------------------------------------------------------------

    DETECT_FIRST_VLAN_TAG_TPID_0 : process(RX_CLIENT_CLK) -- valid by byte 15
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                first_tag_is_vlan_TPID_0_d15   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID0_REG_DATA(16 to 31)) and
                    start_of_frame_array(initial_index + 14) = '1') then
                        first_tag_is_vlan_TPID_0_d15 <= '1';
                    elsif (eof_reset = '1') then
                        first_tag_is_vlan_TPID_0_d15 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a first VLAN tag with type TPID 1
  -------------------------------------------------------------------------

    DETECT_FIRST_VLAN_TAG_TPID_1 : process(RX_CLIENT_CLK) -- valid by byte 15
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                first_tag_is_vlan_TPID_1_d15   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID0_REG_DATA(0 to 15)) and
                    start_of_frame_array(initial_index + 14) = '1') then
                        first_tag_is_vlan_TPID_1_d15 <= '1';
                    elsif (eof_reset = '1') then
                        first_tag_is_vlan_TPID_1_d15 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a first VLAN tag with type TPID 2
  -------------------------------------------------------------------------

    DETECT_FIRST_VLAN_TAG_TPID_2 : process(RX_CLIENT_CLK) -- valid by byte 15
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                first_tag_is_vlan_TPID_2_d15   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID1_REG_DATA(16 to 31)) and
                    start_of_frame_array(initial_index + 14) = '1') then
                        first_tag_is_vlan_TPID_2_d15 <= '1';
                    elsif (eof_reset = '1') then
                        first_tag_is_vlan_TPID_2_d15 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a first VLAN tag with type TPID 3
  -------------------------------------------------------------------------

    DETECT_FIRST_VLAN_TAG_TPID_3 : process(RX_CLIENT_CLK) -- valid by byte 15
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                first_tag_is_vlan_TPID_3_d15   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID1_REG_DATA(0 to 15)) and
                    start_of_frame_array(initial_index + 14) = '1') then
                        first_tag_is_vlan_TPID_3_d15 <= '1';
                    elsif (eof_reset = '1') then
                        first_tag_is_vlan_TPID_3_d15 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a second VLAN tag with type TPID 0
  -------------------------------------------------------------------------

    DETECT_SECOND_VLAN_TAG_TPID_0 : process(RX_CLIENT_CLK) -- valid by byte 19
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                second_tag_is_vlan_TPID_0_d19   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID0_REG_DATA(16 to 31)) and
                    start_of_frame_array(initial_index + 18) = '1') then
                        second_tag_is_vlan_TPID_0_d19 <= '1';
                    elsif (eof_reset = '1') then
                        second_tag_is_vlan_TPID_0_d19 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a second VLAN tag with type TPID 1
  -------------------------------------------------------------------------

    DETECT_SECOND_VLAN_TAG_TPID_1 : process(RX_CLIENT_CLK) -- valid by byte 19
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                second_tag_is_vlan_TPID_1_d19   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID0_REG_DATA(0 to 15)) and
                    start_of_frame_array(initial_index + 18) = '1') then
                        second_tag_is_vlan_TPID_1_d19 <= '1';
                    elsif (eof_reset = '1') then
                        second_tag_is_vlan_TPID_1_d19 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a second VLAN tag with type TPID 2
  -------------------------------------------------------------------------

    DETECT_SECOND_VLAN_TAG_TPID_2 : process(RX_CLIENT_CLK) -- valid by byte 19
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                second_tag_is_vlan_TPID_2_d19   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID1_REG_DATA(16 to 31)) and
                    start_of_frame_array(initial_index + 18) = '1') then
                        second_tag_is_vlan_TPID_2_d19 <= '1';
                    elsif (eof_reset = '1') then
                        second_tag_is_vlan_TPID_2_d19 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- detect if the frame has a second VLAN tag with type TPID 3
  -------------------------------------------------------------------------

    DETECT_SECOND_VLAN_TAG_TPID_3 : process(RX_CLIENT_CLK) -- valid by byte 19
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                second_tag_is_vlan_TPID_3_d19   <= '0';
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (((rx_data_packed_word(23 downto 16) & rx_data_packed_word(31 downto 24)) = RX_CL_CLK_TPID1_REG_DATA(0 to 15)) and
                    start_of_frame_array(initial_index + 18) = '1') then
                        second_tag_is_vlan_TPID_3_d19 <= '1';
                    elsif (eof_reset = '1') then
                        second_tag_is_vlan_TPID_3_d19 <= '0';
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- Initialize the dual port address for the RXD memory
  -------------------------------------------------------------------------
    RXD_ADDR_CNTR: process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                rxd_mem_addr_cntr  <= rxd_mem_empty_mask;
            elsif (rxd_addr_cntr_load = '1') then
                rxd_mem_addr_cntr  <= unsigned(rxd_mem_next_available4write_ptr_cmb);
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (rxd_addr_cntr_en = '1' and rx_data_packed_ready = '1') then
                        rxd_mem_addr_cntr  <= rxd_mem_addr_cntr + 1;
                    end if;
                end if;
            end if;
        end if;
    end process;

  -------------------------------------------------------------------------
  -- Initialize the dual port address for the RXS memory
  -------------------------------------------------------------------------
    RXS_ADDR_CNTR: process (RX_CLIENT_CLK)
    begin
        if rising_edge(RX_CLIENT_CLK) then
            if RESET2RX_CLIENT = '1' then
                rxs_mem_addr_cntr  <= rxs_mem_four_mask;
            elsif (rxs_addr_cntr_load = '1') then
                rxs_mem_addr_cntr  <= unsigned(rxs_mem_next_available4write_ptr_cmb);
            else
                if (RX_CLIENT_CLK_ENBL = '1') then
                    if (rxs_addr_cntr_en = '1' and not(rxs_mem_addr_cntr = rxs_mem_full_mask)) then
                        rxs_mem_addr_cntr  <= rxs_mem_addr_cntr + 1;
                    elsif (rxs_addr_cntr_en = '1' and rxs_mem_addr_cntr = rxs_mem_full_mask) then
                        rxs_mem_addr_cntr  <= rxs_mem_four_mask;
                    end if;
                end if;
            end if;
        end if;
    end process;

    RX_CLIENT_RXS_DPMEM_ADDR(C_RXS_MEM_ADDR_WIDTH downto 0) <=
    std_logic_vector(rxs_mem_one_mask)   when receive_frame_current_state = RESET_INIT_MEM_PTR_2 else
    std_logic_vector(rxs_mem_two_mask)   when receive_frame_current_state = RESET_INIT_MEM_PTR_3 else
    std_logic_vector(rxs_mem_three_mask) when receive_frame_current_state = RESET_INIT_MEM_PTR_4 else
    std_logic_vector(rxs_mem_two_mask)   when receive_frame_current_state = UPDATE_MEM_PTR_2 else
    std_logic_vector(rxs_mem_addr_cntr);

    RX_CLIENT_RXS_DPMEM_WR_EN(0) <=
   '1'  when receive_frame_current_state = RESET_INIT_MEM_PTR_2 else
   '1'  when receive_frame_current_state = RESET_INIT_MEM_PTR_3 else
   '1'  when receive_frame_current_state = RESET_INIT_MEM_PTR_4 else
   '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_1 else
   '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_2 else
   '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_3 else
   '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_4 else
   '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_5 else
   '1'  when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_6 else
   '1'  when receive_frame_current_state = UPDATE_MEM_PTR_2 else
   '0';

   RX_CLIENT_RXS_DPMEM_WR_DATA(35 downto 0) <=
   zero_extend_rxd_mask36 & rxd_mem_last_read_out_ptr_cmb        when receive_frame_current_state = RESET_INIT_MEM_PTR_2 else
   zero_extend_rxs_mask36 & rxs_mem_next_available4write_ptr_cmb when receive_frame_current_state = RESET_INIT_MEM_PTR_3 else
   zero_extend_rxs_mask36 & std_logic_vector(rxs_mem_full_mask)  when receive_frame_current_state = RESET_INIT_MEM_PTR_4 else
   zero_extend_rxs_mask36 & rxs_mem_next_available4write_ptr_cmb when receive_frame_current_state = UPDATE_MEM_PTR_2 else
   rxs_status_word_1_cmb                                         when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_1 else
   rxs_status_word_2                                             when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_2 else
   rxs_status_word_3                                             when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_3 else
   rxs_status_word_4                                             when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_4 else
   rxs_status_word_5                                             when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_5 else
   rxs_status_word_6_cmb                                         when receive_frame_current_state = UPDATE_STATUS_FIFO_WORD_6 else
   (others => '0');

   RX_CLIENT_RXD_DPMEM_WR_EN(0) <=
  rx_data_packed_ready when receive_frame_data_current_state = RECEIVING_FRAME else
  '0';

  RX_CLIENT_RXD_DPMEM_ADDR(C_RXD_MEM_ADDR_WIDTH downto 0) <= std_logic_vector(rxd_mem_addr_cntr);

  RX_CLIENT_RXD_DPMEM_WR_DATA(35 downto 0) <= rx_data_vld_packed_word & rx_data_packed_word;

  --------------------------------------------------------------------------
  -- receive frame State Machine
  -- RXFRMSM_REGS_PROCESS: registered process of the state machine
  -- RXFRMSM_CMB_PROCESS:  combinatorial next-state logic
  --------------------------------------------------------------------------

  RXFRMSM_REGS_PROCESS: process (RX_CLIENT_CLK)
  begin
      if rising_edge(RX_CLIENT_CLK) then
          if RESET2RX_CLIENT = '1' then
              receive_frame_current_state          <= RESET_INIT_MEM_PTR_1;
	      receive_frame_data_current_state     <= RESET;
              rxd_mem_next_available4write_ptr_reg <= std_logic_vector(rxd_mem_empty_mask);
              rxd_mem_last_read_out_ptr_reg        <= std_logic_vector(rxd_mem_full_mask);
              rxs_mem_next_available4write_ptr_reg <= std_logic_vector(rxs_mem_four_mask);
              rxs_status_word_1_reg                <= (others => '0');
              rxs_status_word_6_reg                <= (others => '0');
          else
              if (RX_CLIENT_CLK_ENBL = '1') then
                  receive_frame_current_state          <= receive_frame_next_state;
		  receive_frame_data_current_state     <= receive_frame_data_next_state;
                  rxd_mem_next_available4write_ptr_reg <= rxd_mem_next_available4write_ptr_cmb;
                  rxd_mem_last_read_out_ptr_reg        <= rxd_mem_last_read_out_ptr_cmb;
                  rxs_mem_next_available4write_ptr_reg <= rxs_mem_next_available4write_ptr_cmb;
                  rxs_status_word_1_reg                <= rxs_status_word_1_cmb;
                  rxs_status_word_6_reg                <= rxs_status_word_6_cmb;
              end if;
          end if;
      end if;
  end process;

  RX_RECEIVEFSM_CMD_PROCESS: process (
      receive_frame_data_current_state,  
      rxd_mem_next_available4write_ptr_cmb,
      rxd_mem_next_available4write_ptr_reg,
      rxd_mem_empty_mask,
      rxd_mem_full_mask,
      rxd_mem_last_read_out_ptr_cmb,
      rxd_mem_last_read_out_ptr_reg,
      rxclclk_rxd_mem_last_read_out_ptr_d1,
      rxs_status_word_1_cmb,
      rxs_status_word_1_reg, not_enough_rxs_memory,
      start_of_frame_array,
      end_of_frame_array,
      rxd_mem_addr_cntr,
      save_rx_goodframe,
      save_rx_badframe,
      rx_data_packed_ready,
      rxs_status_word_6_reg,
      RX_CL_CLK_BRDCAST_REJ,
      RX_CL_CLK_MULCAST_REJ,
      frame_is_broadcast_d10,
      frame_is_multicast_d10,
      saveExtendedMulticastReject,
      frame_length_bytes_lat,
      RX_CL_CLK_BAD_FRAME_ENBL
  ) 
  begin
      rxd_addr_cntr_en              <= '0';
      rxd_addr_cntr_load            <= '0';
      RX_FRAME_RECEIVED_INTRPT      <= '0';
      RX_FRAME_REJECTED_INTRPT      <= '0';
      RX_BUFFER_MEM_OVERFLOW_INTRPT <= '0';
      update_status_fifo            <= '0';

      rxd_mem_next_available4write_ptr_cmb <= rxd_mem_next_available4write_ptr_reg;
      rxd_mem_last_read_out_ptr_cmb        <= rxd_mem_last_read_out_ptr_reg;
      rxs_status_word_1_cmb                <= rxs_status_word_1_reg;
      rxs_status_word_6_cmb(15 downto 0)   <= rxs_status_word_6_reg(15 downto 0);
      case receive_frame_data_current_state is
          when RESET =>
              receive_frame_data_next_state        <= WAIT_FOR_START_OF_FRAME;
              rxd_mem_next_available4write_ptr_cmb <= std_logic_vector(rxd_mem_empty_mask);
              rxd_mem_last_read_out_ptr_cmb        <= std_logic_vector(rxd_mem_full_mask);
              rxs_status_word_1_cmb                <= (others => '0');
       
          when WAIT_FOR_START_OF_FRAME =>
              rxd_mem_last_read_out_ptr_cmb    <= rxclclk_rxd_mem_last_read_out_ptr_d1(C_RXD_MEM_ADDR_WIDTH downto 0);
              rxd_addr_cntr_load               <= '1';
              if (start_of_frame_array (1) = '1') then
                  receive_frame_data_next_state    <= RECEIVING_FRAME;
              else
                  receive_frame_data_next_state    <= WAIT_FOR_START_OF_FRAME;
              end if;

          when RECEIVING_FRAME =>
              rxd_mem_last_read_out_ptr_cmb    <= rxclclk_rxd_mem_last_read_out_ptr_d1(C_RXD_MEM_ADDR_WIDTH downto 0);
              rxs_status_word_1_cmb(15 downto C_RXD_MEM_ADDR_WIDTH+1) <= (others => '0');
              rxs_status_word_1_cmb(C_RXD_MEM_ADDR_WIDTH downto 0)    <= rxd_mem_next_available4write_ptr_cmb;
              rxd_addr_cntr_en                 <= '1';
              if (std_logic_vector(rxd_mem_addr_cntr) = rxd_mem_last_read_out_ptr_cmb and rx_data_packed_ready = '1') then -- RXD memory overflow
                  receive_frame_data_next_state    <= WAIT_FOR_START_OF_FRAME;
                  RX_BUFFER_MEM_OVERFLOW_INTRPT  <= '1';
              elsif (end_of_frame_array (1) = '0') then
                  receive_frame_data_next_state    <= RECEIVING_FRAME;
              else
                  receive_frame_data_next_state    <= END_OF_FRAME_CHECK_GOOD_BAD;
              end if;

          when END_OF_FRAME_CHECK_GOOD_BAD =>
              rxs_status_word_1_cmb(35 downto 32)  <= (others => '0');
              rxs_status_word_1_cmb(31 downto 16)  <= std_logic_vector(frame_length_bytes_lat);
              rxs_status_word_6_cmb(15 downto 0)   <= std_logic_vector(frame_length_bytes_lat);
              if (not_enough_rxs_memory = '1') then  -- RXS memory overflow
                  receive_frame_data_next_state    <= WAIT_FOR_START_OF_FRAME;
                  RX_BUFFER_MEM_OVERFLOW_INTRPT  <= '1';
              elsif ((save_rx_goodframe = '1') or (save_rx_badframe = '1' and RX_CL_CLK_BAD_FRAME_ENBL = '1'))  then
                  if ((frame_is_broadcast_d10 = '1' and RX_CL_CLK_BRDCAST_REJ = '1') or
                  (frame_is_multicast_d10 = '1' and RX_CL_CLK_MULCAST_REJ = '1') or
                  (saveExtendedMulticastReject = '1'))then
                      receive_frame_data_next_state       <= WAIT_FOR_START_OF_FRAME;
                      RX_FRAME_REJECTED_INTRPT       <= '1';
                  else
                      rxd_mem_next_available4write_ptr_cmb <= std_logic_vector(rxd_mem_addr_cntr);
                      receive_frame_data_next_state  <= WAIT_FOR_START_OF_FRAME;
                      update_status_fifo             <= '1';
                      RX_FRAME_RECEIVED_INTRPT       <= '1';
                  end if;
              elsif (save_rx_badframe = '1') then
                  receive_frame_data_next_state  <= WAIT_FOR_START_OF_FRAME;
                  RX_FRAME_REJECTED_INTRPT       <= '1';
              else
                  receive_frame_data_next_state  <= END_OF_FRAME_CHECK_GOOD_BAD;
              end if;

      when others   =>
        receive_frame_data_next_state    <= WAIT_FOR_START_OF_FRAME;
      end case;
  end process;

  RXFRMSM_CMB_PROCESS: process (
      receive_frame_current_state,
      rxs_mem_addr_cntr,
      rxs_mem_next_available4write_ptr_cmb, rxs_mem_next_available4write_ptr_reg,
      update_status_fifo,
      rxs_mem_four_mask
  )
  begin

      rxs_addr_cntr_en              <= '0';
      rxs_addr_cntr_load            <= '0';
      rxs_mem_next_available4write_ptr_cmb <= rxs_mem_next_available4write_ptr_reg;


      case receive_frame_current_state is

          when RESET_INIT_MEM_PTR_1 =>
              receive_frame_next_state             <= RESET_INIT_MEM_PTR_2;
              rxs_mem_next_available4write_ptr_cmb <= std_logic_vector(rxs_mem_four_mask);

          when RESET_INIT_MEM_PTR_2 =>
              receive_frame_next_state         <= RESET_INIT_MEM_PTR_3;

          when RESET_INIT_MEM_PTR_3 =>
              receive_frame_next_state         <= RESET_INIT_MEM_PTR_4;

          when RESET_INIT_MEM_PTR_4 =>
              receive_frame_next_state         <= IDLE;

          when IDLE => 
              if (update_status_fifo = '1') then
                  receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_1;
              else
                  receive_frame_next_state         <= IDLE;
              end if;
              rxs_addr_cntr_load               <= '1';

          when UPDATE_STATUS_FIFO_WORD_1 =>
              receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_2;
              rxs_addr_cntr_en                 <= '1';

          when UPDATE_STATUS_FIFO_WORD_2 =>
              receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_3;
              rxs_addr_cntr_en                 <= '1';

          when UPDATE_STATUS_FIFO_WORD_3 =>
              receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_4;
              rxs_addr_cntr_en                 <= '1';

          when UPDATE_STATUS_FIFO_WORD_4 =>
              receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_5;
              rxs_addr_cntr_en                 <= '1';

          when UPDATE_STATUS_FIFO_WORD_5 =>
              receive_frame_next_state         <= UPDATE_STATUS_FIFO_WORD_6;
              rxs_addr_cntr_en                 <= '1';

          when UPDATE_STATUS_FIFO_WORD_6 =>
              receive_frame_next_state         <= UPDATE_MEM_PTR_1;
              rxs_addr_cntr_en                 <= '1';

          when UPDATE_MEM_PTR_1 =>
              receive_frame_next_state         <= UPDATE_MEM_PTR_2;
              rxs_mem_next_available4write_ptr_cmb <= std_logic_vector(rxs_mem_addr_cntr);

          when UPDATE_MEM_PTR_2 =>
              receive_frame_next_state         <= IDLE;

          when others   =>
              receive_frame_next_state         <= RESET_INIT_MEM_PTR_1;
      end case;
  end process;

  -------------------------------------------------------------------------
  -- check enhanced multicast address filtering or not
  -------------------------------------------------------------------------

  EXTENDED_MULTICAST: if(C_MCAST_EXTEND = 1) generate

      type EMCFLTRSM_TYPE is (
      WAIT_FRAME_START,
      GET_SECOND_BYTE,
      GET_THIRD_BYTE,
      GET_FORTH_BYTE,
      GET_FIFTH_BYTE,
      READ_TABLE_ENTRY,
      READ_TABLE_ENTRY2,
      GET_UNI_ADDRESS,
      CHECK_UNI_ADDRESS,
      GET_BRDCAST_ADDRESS,
      CHECK_BRDCAST_ADDRESS,
      ACCEPT_AND_WAIT_TILL_END,
      REJECT_AND_WAIT_TILL_END
  );

  signal eMcFltrSM_Cs           : EMCFLTRSM_TYPE;
  signal eMcFltrSM_Ns           : EMCFLTRSM_TYPE;
  signal tempDestAddr           : std_logic_vector(0 to 47);
  signal unicastMatch           : std_logic;
  signal broadcastMatch         : std_logic;
  signal emacClientRxdLegacy_d1 : std_logic_vector(7 downto 0);

  signal rxClClkMcastEn_i        : std_logic;
  signal rxClClkMcastAddr_i      : std_logic_vector(0 to 14);
  signal rxClClkMcastAddr_i_d    : std_logic_vector(0 to 14);
  signal rx_cl_clk_mcast_rd_data_d1 : std_logic;

  begin

      RX_CL_CLK_MCAST_EN   <= rxClClkMcastEn_i;
      RX_CL_CLK_MCAST_ADDR <= rxClClkMcastAddr_i;

      process(RX_CLIENT_CLK)
      begin
          if(rising_edge(RX_CLIENT_CLK)) then
              if(RESET2RX_CLIENT='1') then
                  emacClientRxdLegacy_d1     <= (others => '0');
                  rx_cl_clk_mcast_rd_data_d1 <= '0';
              else
                  rx_cl_clk_mcast_rd_data_d1 <= RX_CL_CLK_MCAST_RD_DATA(0);
                  if(RX_CLIENT_CLK_ENBL='1') then
                      emacClientRxdLegacy_d1   <= EMAC_CLIENT_RXD_LEGACY;
                  end if;
              end if;
          end if;
      end process;

      COMPARE_UNICAST_ADDR_PROCESS: process (RX_CLIENT_CLK)
      begin
          if (RX_CLIENT_CLK'event and RX_CLIENT_CLK = '1') then
              if (RESET2RX_CLIENT = '1') then
                  unicastMatch <= '0';
              else
                  if (tempDestAddr(0 to 7)   = RX_CL_CLK_UAWL_REG_DATA(24 to 31) and
                  tempDestAddr(8 to 15)  = RX_CL_CLK_UAWL_REG_DATA(16 to 23) and
                  tempDestAddr(16 to 23) = RX_CL_CLK_UAWL_REG_DATA(8 to 15) and
                  tempDestAddr(24 to 31) = RX_CL_CLK_UAWL_REG_DATA(0 to 7) and
                  tempDestAddr(32 to 39) = RX_CL_CLK_UAWU_REG_DATA(24 to 31) and
                  tempDestAddr(40 to 47) = RX_CL_CLK_UAWU_REG_DATA(16 to 23))then
                      unicastMatch <= '1';
                  else
                      unicastMatch <= '0';
                  end if;
              end if;
          end if;
      end process;

      COMPARE_BROADCAST_ADDR_PROCESS: process (RX_CLIENT_CLK)
      begin
          if (RX_CLIENT_CLK'event and RX_CLIENT_CLK = '1') then
              if (RESET2RX_CLIENT = '1') then
                  broadcastMatch <= '0';
              else
                  if (tempDestAddr=x"ffffffffffff") then
                      broadcastMatch <= '1';
                  else
                      broadcastMatch <= '0';
                  end if;
              end if;
          end if;
      end process;

      CAPTURE_TEMPDESTADDR_PROCESS: process (RX_CLIENT_CLK)
      begin
          if (RX_CLIENT_CLK'event and RX_CLIENT_CLK = '1') then
              if (RESET2RX_CLIENT = '1') then
                  tempDestAddr    <= (others => '0');
              else
                  if (RX_CLIENT_CLK_ENBL = '1') then
                      if (start_of_frame_array (initial_index + 1) = '1') then
                          tempDestAddr(0 to 7)   <= emacClientRxdLegacy_d1(7 downto 0);
                          tempDestAddr(8 to 47)  <= (others => '0');
                      elsif (start_of_frame_array (initial_index + 2) = '1') then
                          tempDestAddr(0 to 7)   <= tempDestAddr(0 to 7);
                          tempDestAddr(8 to 15)  <= emacClientRxdLegacy_d1(7 downto 0);
                          tempDestAddr(16 to 47) <= (others => '0');
                      elsif (start_of_frame_array (initial_index + 3) = '1') then
                          tempDestAddr(0 to 15)  <= tempDestAddr(0 to 15);
                          tempDestAddr(16 to 23) <= emacClientRxdLegacy_d1(7 downto 0);
                          tempDestAddr(24 to 47) <= (others => '0');
                      elsif (start_of_frame_array (initial_index + 4) = '1') then
                          tempDestAddr(0 to 23)  <= tempDestAddr(0 to 23);
                          tempDestAddr(24 to 31) <= emacClientRxdLegacy_d1(7 downto 0);
                          tempDestAddr(32 to 47) <= (others => '0');
                      elsif (start_of_frame_array (initial_index + 5) = '1') then
                          tempDestAddr(0 to 31)  <= tempDestAddr(0 to 31);
                          tempDestAddr(32 to 39) <= emacClientRxdLegacy_d1(7 downto 0);
                          tempDestAddr(40 to 47) <= (others => '0');
                      elsif (start_of_frame_array (initial_index + 6) = '1') then
                          tempDestAddr(0 to 39)  <= tempDestAddr(0 to 39);
                          tempDestAddr(40 to 47) <= emacClientRxdLegacy_d1(7 downto 0);
                      else
                          tempDestAddr(0 to 47)  <= tempDestAddr(0 to 47);
                      end if;
                  end if;
              end if;
          end if;
      end process;

  -------------------------------------------------------------------------
  -- save the indication that we had an extended multicast reject
  -------------------------------------------------------------------------

      SAVE_EXTENDED_MULTICAST_REJECT : process(RX_CLIENT_CLK)
      begin
          if rising_edge(RX_CLIENT_CLK) then
              if RESET2RX_CLIENT = '1' then
                  saveExtendedMulticastReject   <= '0';
              else
                  if (eof_reset = '1') then
                      saveExtendedMulticastReject <= '0';
                  elsif (extendedMulticastReject = '1') then
                      saveExtendedMulticastReject <= '1';
                  end if;
              end if;
          end if;
      end process;

      EMCFLTRSM_REGS_PROCESS: process (RX_CLIENT_CLK )
      begin
          if (RX_CLIENT_CLK'event and RX_CLIENT_CLK = '1') then
              if (RESET2RX_CLIENT = '1') then
                  eMcFltrSM_Cs     <= WAIT_FRAME_START;
                  rxClClkMcastAddr_i_d <= (others => '0');
              else
                  if (RX_CLIENT_CLK_ENBL = '1') then
                      eMcFltrSM_Cs <= eMcFltrSM_Ns;
                      rxClClkMcastAddr_i_d <= rxClClkMcastAddr_i;
                  end if;
              end if;
          end if;
      end process;

      EMCFLTRSM_CMB_PROCESS: process (
          eMcFltrSM_Cs,
          start_of_frame_array,
          end_of_frame_array (1),
          RX_CL_CLK_NEW_FNC_ENBL,
          RX_CL_CLK_EMULTI_FLTR_ENBL,
          emacClientRxdLegacy_d1,
          RX_CL_CLK_MCAST_RD_DATA,
          rx_cl_clk_mcast_rd_data_d1,
          tempDestAddr,
          RX_CL_CLK_UAWL_REG_DATA,
          RX_CL_CLK_UAWU_REG_DATA,
          unicastMatch, initial_index,
          rxClClkMcastAddr_i_d,
          rxClClkMcastAddr_i,
          broadcastMatch,
          eof_reset
      )
      begin

          extendedMulticastReject   <= '0';
          rxClClkMcastEn_i          <= '0';
          rxClClkMcastAddr_i        <= rxClClkMcastAddr_i_d;

          case eMcFltrSM_Cs is

              when WAIT_FRAME_START =>
                  rxClClkMcastAddr_i <= (others => '0');
                  if (RX_CL_CLK_NEW_FNC_ENBL = '1' and RX_CL_CLK_EMULTI_FLTR_ENBL = '1') then
                      if (start_of_frame_array (initial_index + 1) = '1')then
                          if (emacClientRxdLegacy_d1=X"01")then
                              eMcFltrSM_Ns <= GET_SECOND_BYTE; -- looks like IP generated multicast so far
                          elsif (emacClientRxdLegacy_d1(0)='0')then
                              eMcFltrSM_Ns <= GET_UNI_ADDRESS; -- it's a unicast address that we need to compare
                          elsif (emacClientRxdLegacy_d1=X"FF")then
                              eMcFltrSM_Ns <= GET_BRDCAST_ADDRESS; -- looks like broadcast so far
                          else
                              eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END; -- must be multicast but non-IP generated
                              extendedMulticastReject <= '1';
                          end if;
                      else
                          eMcFltrSM_Ns <= WAIT_FRAME_START; -- a new frame hasn't started yet
                      end if;
                  else
                      eMcFltrSM_Ns <= WAIT_FRAME_START; -- extended multicast filtering not enabled
                  end if;

              when GET_SECOND_BYTE =>
                  if (emacClientRxdLegacy_d1=X"00")then
                      eMcFltrSM_Ns <= GET_THIRD_BYTE; -- still looks like IP generated multicast so far
                  else
                      eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END; -- must be multicast but non-IP generated
                      extendedMulticastReject <= '1';
                  end if;

              when GET_THIRD_BYTE =>
                  if (emacClientRxdLegacy_d1=X"5e")then
                      eMcFltrSM_Ns <= GET_FORTH_BYTE; -- it is an IP generated multicast so let get the rest and look it up
                  else
                      eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END; -- must be multicast but non-IP generated
                      extendedMulticastReject <= '1';
                  end if;

              when GET_FORTH_BYTE =>
                  rxClClkMcastAddr_i(0 to 6) <= emacClientRxdLegacy_d1(6 downto 0);
                  eMcFltrSM_Ns <= GET_FIFTH_BYTE;

              when GET_FIFTH_BYTE =>
                  rxClClkMcastAddr_i(7 to 14) <= emacClientRxdLegacy_d1(7 downto 0);
                  rxClClkMcastEn_i            <= '1';
                  eMcFltrSM_Ns <= READ_TABLE_ENTRY;

              when READ_TABLE_ENTRY =>
          --rxClClkMcastAddr_i(7 to 14) <= emacClientRxdLegacy_d1(7 downto 0);
                  rxClClkMcastEn_i            <= '1';
                  eMcFltrSM_Ns <= READ_TABLE_ENTRY2;

              when READ_TABLE_ENTRY2 =>
                  rxClClkMcastEn_i            <= '1';
                  if (rx_cl_clk_mcast_rd_data_d1 ='0')then
                      eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END;
                      extendedMulticastReject  <= '1';
                  else
                      eMcFltrSM_Ns <= ACCEPT_AND_WAIT_TILL_END;
                  end if;

              when GET_UNI_ADDRESS =>
                  if (start_of_frame_array (initial_index + 8)='1')then
                      eMcFltrSM_Ns <= CHECK_UNI_ADDRESS;
                  else
                      eMcFltrSM_Ns <= GET_UNI_ADDRESS;
                  end if;

              when GET_BRDCAST_ADDRESS =>
                  if (start_of_frame_array (initial_index + 8)='1')then
                      eMcFltrSM_Ns <= CHECK_BRDCAST_ADDRESS;
                  else
                      eMcFltrSM_Ns <= GET_BRDCAST_ADDRESS;
                  end if;

              when CHECK_BRDCAST_ADDRESS =>
                  if (broadcastMatch='1')then
                      eMcFltrSM_Ns <= ACCEPT_AND_WAIT_TILL_END;
                  else
                      eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END;
                      extendedMulticastReject  <= '1';
                  end if;

              when CHECK_UNI_ADDRESS =>
                  if (unicastMatch = '1')then
                      eMcFltrSM_Ns <= ACCEPT_AND_WAIT_TILL_END;
                  else
                      eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END;
                      extendedMulticastReject  <= '1';
                  end if;

              when REJECT_AND_WAIT_TILL_END =>
                  if (eof_reset = '1' )then
                      eMcFltrSM_Ns <= WAIT_FRAME_START;
                      extendedMulticastReject  <= '0';
                  else
                      eMcFltrSM_Ns <= REJECT_AND_WAIT_TILL_END;
                      extendedMulticastReject  <= '1';
                  end if;

              when ACCEPT_AND_WAIT_TILL_END =>
                  extendedMulticastReject  <= '0';
                  if (eof_reset = '1' )then
                      eMcFltrSM_Ns <= WAIT_FRAME_START;
                  else
                      eMcFltrSM_Ns <= ACCEPT_AND_WAIT_TILL_END;
                  end if;

              when others   =>
                  eMcFltrSM_Ns <= WAIT_FRAME_START;
          end case;
      end process;


  end generate EXTENDED_MULTICAST;

  NO_EXTENDED_MULTICAST: if(C_MCAST_EXTEND = 0) generate
  begin
      extendedMulticastReject <= '0';
      RX_CL_CLK_MCAST_ADDR    <= (others => '0');
      RX_CL_CLK_MCAST_EN      <= '0';
      saveExtendedMulticastReject   <= '0';
  end generate NO_EXTENDED_MULTICAST;

end rtl;



------------------------------------------------------------------------------
-- rx_axistream_if.vhd
------------------------------------------------------------------------------
-- (c) Copyright 2004-2009 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, rtlLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-- ------------------------------------------------------------------------------
--
------------------------------------------------------------------------------
-- Filename:        rx_axistream_if.vhd
-- Version:         v1.00a
-- Description:     Receive interface between AXIStream and Temac
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to rtlrove
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:          MSH
--
--  MSH     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of : out   std_logic; port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Libraries used;
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

---library lib_fifo_v1_0;
---use lib_fifo_v1_0.all;
---

library work;
use work.rx_if_pack.all;

-------------------------------------------------------------------------------
-- Definition of Generics :
-------------------------------------------------------------------------------
-- System generics
--  C_FAMILY              -- Xilinx FPGA Family
--  C_RXD_MEM_BYTES               -- Depth of RX memory in Bytes
--  C_RXCSUM
--     0  No checksum offloading
--     1  Partial (legacy) checksum offloading
--     2  Full checksum offloading
--  C_RXVLAN_TRAN         -- Enable RX enhanced VLAN translation
--  C_RXVLAN_TAG          -- Enable RX enhanced VLAN taging
--  C_RXVLAN_STRP         -- Enable RX enhanced VLAN striping
--  C_MCAST_EXTEND        -- Enable RX extended multicast address filtering

-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Definition of Ports :
-------------------------------------------------------------------------------
--    BUS2IP_CLK
--    BUS2IP_RESET
--
--    AXI_STR_RXD_ACLK
--    AXI_STR_RXD_VALID
--    AXI_STR_RXD_READY
--    AXI_STR_RXD_LAST
--    AXI_STR_RXD_STRB
--    AXI_STR_RXD_DATA
--
--    AXI_STR_RXS_ACLK
--    AXI_STR_RXS_VALID
--    AXI_STR_RXS_READY
--    AXI_STR_RXS_LAST
--    AXI_STR_RXS_STRB
--    AXI_STR_RXS_DATA
--
--    EMAC_CLIENT_RXD_LEGACY
--    EMAC_CLIENT_RXD_VLD_LEGACY
--    EMAC_CLIENT_RX_GOODFRAME_LEGACY
--    EMAC_CLIENT_RX_BADFRAME_LEGACY
--    EMAC_CLIENT_RX_FRAMEDROP
--    LEGACY_RX_FILTER_MATCH
--
--    RX_CLIENT_CLK
--    RX_CLIENT_CLK_ENBL
--
--    EMAC_CLIENT_RX_STATS
--    EMAC_CLIENT_RX_STATS_VLD
--    EMAC_CLIENT_RX_STATS_BYTE_VLD
--    EMAC_CLIENT_RXD_VLD_2STATS
--    SOFT_EMAC_CLIENT_RX_STATS
--
--    RTAGREGDATA
--    TPID0REGDATA
--    TPID1REGDATA
--    UAWLREGDATA
--    UAWUREGDATA
--    RXCLCLKMCASTADDR
--    RXCLCLKMCASTEN
--    RXCLCLKMCASTRDDATA
--    LLINKCLKVLANADDR
--    LLINKCLKVLANRDDATA
--    LLINKCLKRXVLANBRAMENA
--
--    LLINKCLKEMULTIFLTRENBL
--    LLINKCLKNEWFNCENBL
--    LLINKCLKRXVSTRPMODE
--    LLINKCLKRXVTAGMODE
-------------------------------------------------------------------------------
----                  Entity Section
-------------------------------------------------------------------------------

entity rx_axistream_if is
  generic (
    C_RXD_MEM_BYTES       : integer                       := 4096;
    C_RXD_MEM_ADDR_WIDTH  : integer                       := 10;
    C_RXS_MEM_BYTES       : integer                       := 4096;
    C_RXS_MEM_ADDR_WIDTH  : integer                       := 10;
    C_FAMILY              : string                        := "virtex6";
    C_RXCSUM              : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_RXVLAN_TRAN         : integer range 0 to 1          := 0;
    C_RXVLAN_TAG          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP         : integer range 0 to 1          := 0;
    C_MCAST_EXTEND        : integer range 0 to 1          := 0
    );

  port    (
    AXI_STR_RXD_ACLK                : in  std_logic;                                        --  Receive AXI-Stream Data Clock
    AXI_STR_RXD_VALID               : out std_logic;                                        --  Receive AXI-Stream Data VALID
    AXI_STR_RXD_READY               : in  std_logic;                                        --  Receive AXI-Stream Data READY
    AXI_STR_RXD_LAST                : out std_logic;                                        --  Receive AXI-Stream Data LAST
    AXI_STR_RXD_STRB                : out std_logic_vector(3 downto 0);                     --  Receive AXI-Stream Data STRB
    AXI_STR_RXD_DATA                : out std_logic_vector(31 downto 0);                    --  Receive AXI-Stream Data DATA
    RESET2AXI_STR_RXD               : in  std_logic;                                        --  Reset

    AXI_STR_RXS_ACLK                : in  std_logic;                                        --  Receive AXI-Stream Status Clock
    AXI_STR_RXS_VALID               : out std_logic;                                        --  Receive AXI-Stream Status VALID
    AXI_STR_RXS_READY               : in  std_logic;                                        --  Receive AXI-Stream Status READY
    AXI_STR_RXS_LAST                : out std_logic;                                        --  Receive AXI-Stream Status LAST
    AXI_STR_RXS_STRB                : out std_logic_vector(3 downto 0);                     --  Receive AXI-Stream Status STRB
    AXI_STR_RXS_DATA                : out std_logic_vector(31 downto 0);                    --  Receive AXI-Stream Status DATA
    RESET2AXI_STR_RXS               : in  std_logic;                                        --  Reset

    AXI_STR_RXD_DPMEM_WR_DATA       : out std_logic_vector(35 downto 0);                    --  Receive Data Memory Wr Data
    AXI_STR_RXD_DPMEM_RD_DATA       : in  std_logic_vector(35 downto 0);                    --  Receive Data Memory Rd Data
    AXI_STR_RXD_DPMEM_WR_EN         : out std_logic_vector(0 downto 0);                     --  Receive Data Memory Wr Enable
    AXI_STR_RXD_DPMEM_ADDR          : out std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  Receive Data Memory Addr

    AXI_STR_RXS_DPMEM_WR_DATA       : out std_logic_vector(35 downto 0);                    --  Receive Status Memory Wr Data
    AXI_STR_RXS_DPMEM_RD_DATA       : in  std_logic_vector(35 downto 0);                    --  Receive Status Memory Rd Data
    AXI_STR_RXS_DPMEM_WR_EN         : out std_logic_vector(0 downto 0);                     --  Receive Status Memory Wr Enable
    AXI_STR_RXS_DPMEM_ADDR          : out std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  Receive Status Memory Addr

    AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY : out std_logic_vector(35 downto 0);             --  Receive Status GRAY Pointer

	-- The following output is flawed in that the binary version can change by more than 1 value per clock cycle, which means the gray code CDC breaks down.
    AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY : out std_logic_vector(35 downto 0)              --  Receive Data GRAY Pointer
    );
end rx_axistream_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of rx_axistream_if is

---------------------------------------------------------------------
-- Functions
---------------------------------------------------------------------

-- Convert a binary value into a gray code
function bin_to_gray (
   bin : std_logic_vector)
   return std_logic_vector is

   variable gray : std_logic_vector(bin'range);

begin

   for i in bin'range loop
      if i = bin'left then
         gray(i) := bin(i);
      else
         gray(i) := bin(i+1) xor bin(i);
      end if;
   end loop;  -- i

   return gray;

end bin_to_gray;

constant PRE_GRAY_CODED_FF : std_logic_vector(35 downto 0) := x"FFFFFFFFF";

component  basic_sfifo_fg 
  generic (
    C_DWIDTH                      : Integer :=  32 ;
    C_DEPTH                       : Integer := 512 ;
    C_HAS_DATA_COUNT              : integer :=   1 ;
    C_DATA_COUNT_WIDTH            : integer :=  10 ;
    C_IMPLEMENTATION_TYPE         : integer range 0 to 1 := 0;  
    C_MEMORY_TYPE                 : integer := 1;
    C_PRELOAD_REGS                : integer := 1; 
    C_PRELOAD_LATENCY             : integer := 0;              
    C_USE_FWFT_DATA_COUNT         : integer := 0; 
    C_SYNCHRONIZER_STAGE          : integer := 2;   -- valid values are 0 to 8;
    C_FAMILY                      : string  := "virtex6"
    );
  port (
    CLK                           : IN  std_logic := '0';
    DIN                           : IN  std_logic_vector(C_DWIDTH-1 DOWNTO 0) := (OTHERS => '0');
    RD_EN                         : IN  std_logic := '0';  
    SRST                          : IN  std_logic := '0';
    WR_EN                         : IN  std_logic := '0';
    DATA_COUNT                    : OUT std_logic_vector(C_DATA_COUNT_WIDTH-1 DOWNTO 0);
    DOUT                          : OUT std_logic_vector(C_DWIDTH-1 DOWNTO 0);
    EMPTY                         : OUT std_logic;
    FULL                          : OUT std_logic
    );
end component  ;

type RXS_AXISTREAM_STATES is (
  RESET_INIT_1,
  RESET_INIT_2,
  READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_1,
  READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_2,
  ADDR_SETUP_PAUSE_1,
  READ_RXD_MEM_LAST_READ_OUT_PTR,
  ADDR_SETUP_PAUSE_2,
  READ_RXS_MEM_NEXT_AVAILABLE4WRITE_PTR_1,
  READ_RXS_MEM_NEXT_AVAILABLE4WRITE_PTR_2,
  ADDR_SETUP_PAUSE_3,
  READ_RXS_MEM_LAST_READ_OUT_PTR,
  PAUSE_READ_STATUS_WORD1,
  READ_STATUS_WORD1,
  READ_STATUS_WORD2,
  READ_STATUS_WORD3,
  READ_STATUS_WORD4,
  READ_STATUS_WORD5,
  READ_STATUS_WORD6,
  UPDATE_RXS_MEM_LAST_READ_OUT_PTR,
  SEND_STATUS_WORD1,
  SEND_STATUS_WORD2,
  SEND_STATUS_WORD3,
  SEND_STATUS_WORD4,
  SEND_STATUS_WORD5,
  SEND_STATUS_WORD6,
  WAIT_FRAME_DONE,
  UPDATE_RXD_MEM_LAST_READ_OUT_PTR,
  REPEAT_AGAIN
  );

signal rxs_axistream_current_state : RXS_AXISTREAM_STATES;
signal rxs_axistream_next_state    : RXS_AXISTREAM_STATES;

type RXD_AXISTREAM_STATES is (
  IDLE,
  PRIME,
  WRITE_FIRST_WORD,
  LOAD_FIRST_WORD,
  RD_FRAME_FROM_MEM,
  ALMOST_FULL_WAIT1,
  ALMOST_FULL_WAIT2,
  ALMOST_FULL_WAIT3,
  ALMOST_FULL_WAIT4,
  WAIT_END_FRAME,
  PRE_IDLE);

signal rxd_axistream_current_state : RXD_AXISTREAM_STATES;
signal rxd_axistream_next_state    : RXD_AXISTREAM_STATES;

signal rxs_mem_next_available4write_ptr_1_reg : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_next_available4write_ptr_1_cmb : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);

signal rxd_mem_next_available4write_ptr_1_reg : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_next_available4write_ptr_1_cmb : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);

signal axi_str_rxs_dpmem_rd_data_d1           : std_logic_vector(35 downto 0);

signal rxd2rxs_frame_done                     : std_logic;
signal rxs2rxd_frame_done                     : std_logic;

signal frame_length_bytes               : std_logic_vector(15 downto 0);
signal frame_length_words               : integer range 0 to 32767;
signal last_rxd_strb                    : std_logic_vector(3 downto 0);

signal rxd_mem_next_available4write_ptr_cmb : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_next_available4write_ptr_reg : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_last_read_out_ptr_cmb        : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_last_read_out_ptr_reg        : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_next_available4write_ptr_cmb : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_next_available4write_ptr_reg : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_last_read_out_ptr_true_cmb   : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_last_read_out_ptr_true_reg   : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_last_read_out_ptr_cmb        : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_last_read_out_ptr_reg        : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_last_read_out_ptr_plus_one   : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);

signal rxd_mem_full_mask                : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_full_mask_minus_one      : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_empty_mask               : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_one_mask                 : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxd_mem_two_mask                 : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_full_mask                : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_full_mask_minus_one      : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_empty_mask               : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_one_mask                 : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_two_mask                 : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_three_mask               : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_four_mask                : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);

signal zero_extend_rxd_mask36           : std_logic_vector(35 downto C_RXD_MEM_ADDR_WIDTH + 1);
signal zero_extend_rxs_mask36           : std_logic_vector(35 downto C_RXS_MEM_ADDR_WIDTH + 1);

signal rxs_status_word_1                : std_logic_vector(35 downto 0);
signal rxs_status_word_2                : std_logic_vector(35 downto 0);
signal rxs_status_word_3                : std_logic_vector(35 downto 0);
signal rxs_status_word_4                : std_logic_vector(35 downto 0);
signal rxs_status_word_5                : std_logic_vector(35 downto 0);
signal rxs_status_word_6                : std_logic_vector(35 downto 0);

signal rxd_addr_cntr_en                 : std_logic;
signal rxd_mem_addr_cntr                : unsigned(C_RXD_MEM_ADDR_WIDTH downto 0);

signal rxs2rxd_frame_ready              : std_logic;

signal fifoDataIn    : std_logic_vector(0 to 35);
signal fifoWrEn      : std_logic;
signal fifoRdEn      : std_logic;
signal fifoDataOut   : std_logic_vector(0 to 35);
signal fifoDataOut_1d : std_logic_vector(0 to 35) := (others => '0');
signal fifoFull      : std_logic;
signal fifoEmpty     : std_logic;
signal fifoEmpty_1d  : std_logic := '0';
signal fifoDataCount      : std_logic_vector(0 to 5);
signal fifoAlmostFull     : std_logic;
signal rxd_addr_cntr_load : std_logic;
signal rxd_word_cnt       : integer range 0 to 32767;
signal rxd_word_cnt_vector : std_logic_vector (15 downto 0);
signal AXI_STR_RXD_LAST_INT      : std_logic;
signal AXI_STR_RXD_LAST_INT_1D   : std_logic := '0';
signal AXI_STR_RXD_LAST_FED      : std_logic;
signal AXI_STR_RXD_READY_1D      : std_logic := '0';
signal AXI_STR_RXD_READY_RED     : std_logic;
signal LAST_READY_DEASSERT       : std_logic;
signal LAST_READY_DEASSERT_LATCH : std_logic := '0';
signal AXI_STR_RXD_LAST_FALL_LATCH : std_logic := '0';
signal AXI_STR_RXD_STRB_CHK        : std_logic := '0';

signal rxd_mem_last_read_out_ptr_gray_d1           : std_logic_vector(35 downto 0);
signal rxd_mem_last_read_out_ptr_gray              : std_logic_vector(35 downto 0);
signal rxd_mem_last_read_out_ptr_toconvertto_gray  : std_logic_vector(35 downto 0);

signal rxs_mem_last_read_out_ptr_toconvertto_gray        : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_last_read_out_ptr_toconvertto_gray_clean  : unsigned(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_last_read_out_ptr_gray                    : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rxs_mem_last_read_out_ptr_gray_d1                 : std_logic_vector(35 downto 0);

--------------------------------------------------------
-- Declare general attributes used in this file
-- for defining each component being used with
-- the generatecore utility

attribute box_type: string;
attribute GENERATOR_DEFAULT: string;

  -----------------------------------------------------------------------------
  -- The following is the location of the DualPort Memory pointers in the RXS
  -- memory
  -- Address:  Pointer:
  --   0x0       rxd_mem_next_available4write_ptr
  --   0x1       rxd_mem_last_read_out_ptr
  --   0x2       rxs_mem_next_available4write_ptr
  --   0x3       rxs_mem_last_read_out_ptr
  -----------------------------------------------------------------------------


begin

  -------------------------------------------------------------------------
  -- Convert binary encoded RXS last read pointer to gray encoded to send
  -- to receive client interface
  -------------------------------------------------------------------------
  GET_RXS_LAST_READ_GRAY_PROCESS: process (AXI_STR_RXS_ACLK)
  begin
    if rising_edge(AXI_STR_RXS_ACLK) then
      if RESET2AXI_STR_RXS = '1' then
        rxs_mem_last_read_out_ptr_toconvertto_gray <= (others => '0');
      else
        if (rxs_axistream_current_state = READ_STATUS_WORD6 or
            rxs_axistream_current_state = READ_STATUS_WORD1 or
            rxs_axistream_current_state = READ_STATUS_WORD2 or
            rxs_axistream_current_state = READ_STATUS_WORD3 or
            rxs_axistream_current_state = READ_STATUS_WORD4 or
            rxs_axistream_current_state = READ_STATUS_WORD5
        ) then
          rxs_mem_last_read_out_ptr_toconvertto_gray <= rxs_mem_last_read_out_ptr_reg;
        end if;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------------
  -- This processes ensures that the grey code is clean
  -------------------------------------------------------------------------------
  process(AXI_STR_RXS_ACLK)
    begin
      if rising_edge(AXI_STR_RXS_ACLK) then
        if RESET2AXI_STR_RXS = '1' then
          rxs_mem_last_read_out_ptr_toconvertto_gray_clean <= (others => '0');
        else
          if(to_integer(unsigned(rxs_mem_last_read_out_ptr_toconvertto_gray)) > 0) then
            if(rxs_mem_last_read_out_ptr_toconvertto_gray_clean < unsigned(rxs_mem_last_read_out_ptr_toconvertto_gray)) then
              rxs_mem_last_read_out_ptr_toconvertto_gray_clean <= rxs_mem_last_read_out_ptr_toconvertto_gray_clean + 1;
            elsif(rxs_mem_last_read_out_ptr_toconvertto_gray_clean > unsigned(rxs_mem_last_read_out_ptr_toconvertto_gray)) then
              rxs_mem_last_read_out_ptr_toconvertto_gray_clean <= rxs_mem_last_read_out_ptr_toconvertto_gray_clean + 1;
            end if;
        end if;
        end if;
      end if;
  end process;

  rxs_mem_last_read_out_ptr_gray <= bin_to_gray(std_logic_vector(rxs_mem_last_read_out_ptr_toconvertto_gray_clean));

  -------------------------------------------------------------------------
  -- Register gray encoded RXS last read pointer to send to receive client
  -- interface. reset to all ones at power-up
  -------------------------------------------------------------------------
  RXS_LAST_READ_GRAY_PROCESS: process (AXI_STR_RXS_ACLK)
  begin
    if rising_edge(AXI_STR_RXS_ACLK) then
      if RESET2AXI_STR_RXS = '1' then
        rxs_mem_last_read_out_ptr_gray_d1  <= bin_to_gray(PRE_GRAY_CODED_FF);
      else
        rxs_mem_last_read_out_ptr_gray_d1(35 downto C_RXS_MEM_ADDR_WIDTH + 1) <= (others => '0');
        rxs_mem_last_read_out_ptr_gray_d1(C_RXS_MEM_ADDR_WIDTH downto 0) <= rxs_mem_last_read_out_ptr_gray;
      end if;
    end if;
  end process;

  AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY <= rxs_mem_last_read_out_ptr_gray_d1;

  -------------------------------------------------------------------------
  -- Convert binary encoded RXD last read pointer to gray encoded to send
  -- to receive client interface
  -------------------------------------------------------------------------
  rxd_mem_last_read_out_ptr_toconvertto_gray(35 downto C_RXD_MEM_ADDR_WIDTH + 1) <= (others => '0');
  rxd_mem_last_read_out_ptr_toconvertto_gray(C_RXD_MEM_ADDR_WIDTH downto 0) <= std_logic_vector(rxd_mem_addr_cntr - 1) when
    not(rxs_axistream_current_state = UPDATE_RXD_MEM_LAST_READ_OUT_PTR) else
    std_logic_vector(unsigned(rxd_mem_last_read_out_ptr_reg) - 1);
  rxd_mem_last_read_out_ptr_gray <= bin_to_gray(rxd_mem_last_read_out_ptr_toconvertto_gray);

  -------------------------------------------------------------------------
  -- Register gray encoded RXD last read pointer to send to receive client
  -- interface. reset to all ones at power-up
  -------------------------------------------------------------------------
  RXD_LAST_READ_GRAY_PROCESS: process (AXI_STR_RXS_ACLK)
  begin
    if rising_edge(AXI_STR_RXS_ACLK) then
      if RESET2AXI_STR_RXS = '1' then
        rxd_mem_last_read_out_ptr_gray_d1  <= bin_to_gray(PRE_GRAY_CODED_FF);
      else
        if (rxs_axistream_current_state = SEND_STATUS_WORD1 or
            rxs_axistream_current_state = SEND_STATUS_WORD2 or
            rxs_axistream_current_state = SEND_STATUS_WORD3 or
            rxs_axistream_current_state = SEND_STATUS_WORD4 or
            rxs_axistream_current_state = SEND_STATUS_WORD5 or
            rxs_axistream_current_state = SEND_STATUS_WORD6 or
            ((rxs_axistream_current_state = WAIT_FRAME_DONE) and (rxd_addr_cntr_en = '1'))   or
            rxs_axistream_current_state = UPDATE_RXD_MEM_LAST_READ_OUT_PTR
        ) then
          rxd_mem_last_read_out_ptr_gray_d1 <= rxd_mem_last_read_out_ptr_gray;
        end if;
      end if;
    end if;
  end process;

  AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY <= rxd_mem_last_read_out_ptr_gray_d1;

-------------------------------------------------------------------------------

  PIPE_RXS_READ_DATA: process (AXI_STR_RXS_ACLK) -- clock to out of BRAM is slow so register it to make timing easier
  begin
    if rising_edge(AXI_STR_RXS_ACLK) then
      if RESET2AXI_STR_RXS = '1' then
        axi_str_rxs_dpmem_rd_data_d1 <= (others => '0');
      else
        axi_str_rxs_dpmem_rd_data_d1 <= AXI_STR_RXS_DPMEM_RD_DATA;
      end if;
    end if;
  end process;

  -------------------------------------------------------------------------
  -- Generate variable width address masks for checking memory pointers
  -------------------------------------------------------------------------
  RXD_GEN_MASK: for I in C_RXD_MEM_ADDR_WIDTH downto 0 generate
    rxd_mem_full_mask(I) <= '1';
    rxd_mem_empty_mask(I)  <= '0';
  end generate;

  rxd_mem_one_mask            <= rxd_mem_empty_mask + 1;
  rxd_mem_two_mask            <= rxd_mem_empty_mask + 2;
  rxd_mem_full_mask_minus_one <= rxd_mem_full_mask - 1;

  RXS_GEN_MASK: for I in C_RXS_MEM_ADDR_WIDTH downto 0 generate
    rxs_mem_full_mask(I) <= '1';
    rxs_mem_empty_mask(I)  <= '0';
  end generate;

  rxs_mem_one_mask            <= rxs_mem_empty_mask + 1;
  rxs_mem_two_mask            <= rxs_mem_empty_mask + 2;
  rxs_mem_three_mask          <= rxs_mem_empty_mask + 3;
  rxs_mem_four_mask           <= rxs_mem_empty_mask + 4;
  rxs_mem_full_mask_minus_one <= rxs_mem_full_mask - 1;

  zero_extend_rxd_mask36      <= (others => '0');
  zero_extend_rxs_mask36      <= (others => '0');


  RXD_MEM_ADDR_COUNTER: process (AXI_STR_RXD_ACLK)
  begin
    if rising_edge(AXI_STR_RXD_ACLK) then
      if RESET2AXI_STR_RXD = '1' then
        rxd_mem_addr_cntr    <= (others => '0');
      elsif (rxd_addr_cntr_load = '1') then
        rxd_mem_addr_cntr  <= unsigned(rxs_status_word_1(C_RXD_MEM_ADDR_WIDTH downto 0));
      else
        if (rxd_addr_cntr_en = '1') then
          rxd_mem_addr_cntr  <= rxd_mem_addr_cntr + 1;
        end if;
      end if;
    end if;
  end process;

  rxd_word_cnt_vector(15 downto 0) <= std_logic_vector(to_unsigned(rxd_word_cnt,16));

  STORE_STATUS_WORDS: process (AXI_STR_RXS_ACLK)
  --  There is no chance of a simultaneous RXD DPMEM write/read here because at this point this
  --  area of memory has long since been written
  begin
    if rising_edge(AXI_STR_RXS_ACLK) then
      if RESET2AXI_STR_RXS = '1' then
        rxs_status_word_1         <= (others => '0');
        rxs_status_word_2         <= (others => '0');
        rxs_status_word_3         <= (others => '0');
        rxs_status_word_4         <= (others => '0');
        rxs_status_word_5         <= (others => '0');
        rxs_status_word_6         <= (others => '0');
        frame_length_bytes        <= (others => '0');
        frame_length_words        <= 0;
        last_rxd_strb             <= (others => '1');
      else
        if (rxs_axistream_current_state = READ_STATUS_WORD1) then
          rxs_status_word_1  <= axi_str_rxs_dpmem_rd_data_d1;
          frame_length_bytes <= axi_str_rxs_dpmem_rd_data_d1(31 downto 16);
          case axi_str_rxs_dpmem_rd_data_d1(17 downto 16) is
            when "00" =>
              frame_length_words  <= to_integer(unsigned(axi_str_rxs_dpmem_rd_data_d1(31 downto 18)));
              last_rxd_strb       <= x"f";
            when "01" =>
              frame_length_words  <= to_integer(unsigned(axi_str_rxs_dpmem_rd_data_d1(31 downto 18))) + 1;
              last_rxd_strb       <= x"1";
            when "10" =>
              frame_length_words  <= to_integer(unsigned(axi_str_rxs_dpmem_rd_data_d1(31 downto 18))) + 1;
              last_rxd_strb       <= x"3";
            when "11" =>
              frame_length_words  <= to_integer(unsigned(axi_str_rxs_dpmem_rd_data_d1(31 downto 18))) + 1;
              last_rxd_strb       <= x"7";
            -- coverage off
            when others => null;
            -- coverage on
          end case;
        end if;
        if (rxs_axistream_current_state = READ_STATUS_WORD2) then
          rxs_status_word_2  <= AXI_STR_RXS_DPMEM_RD_DATA;
        end if;
        if (rxs_axistream_current_state = READ_STATUS_WORD3) then
          rxs_status_word_3  <= AXI_STR_RXS_DPMEM_RD_DATA;
        end if;
        if (rxs_axistream_current_state = READ_STATUS_WORD4) then
          rxs_status_word_4  <= AXI_STR_RXS_DPMEM_RD_DATA;
        end if;
        if (rxs_axistream_current_state = READ_STATUS_WORD5) then
          rxs_status_word_5  <= AXI_STR_RXS_DPMEM_RD_DATA;
        end if;
        if (rxs_axistream_current_state = READ_STATUS_WORD6) then
          rxs_status_word_6  <= AXI_STR_RXS_DPMEM_RD_DATA;
        end if;
      end if;
    end if;
  end process;

  INC_RXS_MEM_LAST_READ_OUT: process (AXI_STR_RXS_ACLK)
  begin
    if rising_edge(AXI_STR_RXS_ACLK) then
      if RESET2AXI_STR_RXS = '1' then
        rxs_mem_last_read_out_ptr_plus_one <= (others => '1');
      else
        if (rxs_mem_last_read_out_ptr_cmb = rxs_mem_full_mask)then
          rxs_mem_last_read_out_ptr_plus_one <= rxs_mem_four_mask;
        else
          rxs_mem_last_read_out_ptr_plus_one <= rxs_mem_last_read_out_ptr_cmb + 1;
        end if;
      end if;
    end if;
  end process;

  --------------------------------------------------------------------------
  -- receive status AXIStream State Machine
  -- RXSTSSM_REGS_PROCESS: registered process of the state machine
  -- RXSTSSM_CMB_PROCESS:  combinatorial next-state logic
  --------------------------------------------------------------------------

  RXSTSSM_REGS_PROCESS: process (AXI_STR_RXS_ACLK)
  begin
    if rising_edge(AXI_STR_RXS_ACLK) then
      if RESET2AXI_STR_RXS = '1' then
        rxs_axistream_current_state            <= RESET_INIT_1;
        rxd_mem_last_read_out_ptr_reg          <= (others => '0');
        rxs_mem_last_read_out_ptr_reg          <= (others => '0');
        rxs_mem_last_read_out_ptr_true_reg     <= (others => '0');
        rxd_mem_next_available4write_ptr_reg   <= (others => '0');
        rxs_mem_next_available4write_ptr_reg   <= (others => '0');
        rxs_mem_next_available4write_ptr_1_reg <= (others => '0');
        rxd_mem_next_available4write_ptr_1_reg <= (others => '0');
      else
        rxs_axistream_current_state            <= rxs_axistream_next_state;
        rxd_mem_last_read_out_ptr_reg          <= rxd_mem_last_read_out_ptr_cmb;
        rxs_mem_last_read_out_ptr_reg          <= std_logic_vector(rxs_mem_last_read_out_ptr_cmb);
        rxs_mem_last_read_out_ptr_true_reg     <= rxs_mem_last_read_out_ptr_true_cmb;
        rxs_mem_next_available4write_ptr_reg   <= rxs_mem_next_available4write_ptr_cmb;
        rxd_mem_next_available4write_ptr_reg   <= rxd_mem_next_available4write_ptr_cmb;
        rxs_mem_next_available4write_ptr_1_reg <= rxs_mem_next_available4write_ptr_1_cmb;
        rxd_mem_next_available4write_ptr_1_reg <= rxd_mem_next_available4write_ptr_1_cmb;
      end if;
    end if;
  end process;

  RXSTSSM_CMB_PROCESS: process (
    rxs_axistream_current_state,
    AXI_STR_RXS_DPMEM_RD_DATA,
    rxd2rxs_frame_done,
    AXI_STR_RXS_READY,
    rxs_mem_last_read_out_ptr_reg,
    rxs_mem_last_read_out_ptr_cmb,
    rxs_mem_last_read_out_ptr_true_reg,
    rxs_mem_last_read_out_ptr_true_cmb,
    rxd_mem_last_read_out_ptr_reg,
    rxd_mem_last_read_out_ptr_cmb,
    rxs_mem_next_available4write_ptr_reg,
    rxs_mem_next_available4write_ptr_cmb,
    rxd_mem_next_available4write_ptr_reg,
    rxd_mem_next_available4write_ptr_cmb,
    rxs_mem_empty_mask,
    rxs_mem_three_mask,
    rxs_mem_full_mask,
    rxd_addr_cntr_en,
    rxd_mem_addr_cntr,
    rxs_mem_two_mask,
    rxs_mem_one_mask,
    rxs_mem_four_mask,
    rxs_mem_last_read_out_ptr_plus_one,
    rxs_status_word_2,
    rxs_status_word_3,
    rxs_status_word_4,
    rxs_status_word_5,
    rxs_status_word_6,
    axi_str_rxs_dpmem_rd_data_d1,
    rxs_mem_next_available4write_ptr_1_reg,
    rxd_mem_next_available4write_ptr_1_reg,
    rxs_mem_next_available4write_ptr_1_cmb,
    rxd_mem_next_available4write_ptr_1_cmb
    )
  begin
    rxs_mem_last_read_out_ptr_cmb        <= unsigned(rxs_mem_last_read_out_ptr_reg);
    rxd_mem_last_read_out_ptr_cmb        <= rxd_mem_last_read_out_ptr_reg;
    rxs_mem_last_read_out_ptr_true_cmb   <= rxs_mem_last_read_out_ptr_true_reg;
    rxs_mem_next_available4write_ptr_cmb <= rxs_mem_next_available4write_ptr_reg;
    rxd_mem_next_available4write_ptr_cmb <= rxd_mem_next_available4write_ptr_reg;

    rxs_mem_next_available4write_ptr_1_cmb <= rxs_mem_next_available4write_ptr_1_reg;
    rxd_mem_next_available4write_ptr_1_cmb <= rxd_mem_next_available4write_ptr_1_reg;

    AXI_STR_RXD_DPMEM_WR_DATA            <= (others => '0');
    AXI_STR_RXD_DPMEM_WR_EN              <= (others => '0');
    AXI_STR_RXS_DPMEM_WR_DATA            <= (others => '0');
    AXI_STR_RXS_DPMEM_WR_EN              <= (others => '0');
    AXI_STR_RXS_DPMEM_ADDR               <= std_logic_vector(rxs_mem_three_mask); -- rxs_mem_last_read_out_ptr
    rxs2rxd_frame_ready                  <= '0';
    AXI_STR_RXS_VALID                    <= '0';
    AXI_STR_RXS_LAST                     <= '0';
    AXI_STR_RXS_STRB                     <= X"F";
    AXI_STR_RXS_DATA                     <= (others => '0');

    case rxs_axistream_current_state is

      when RESET_INIT_1 =>
      -- we must wait until the rx client interface has initialized the ptrs in dpmem;
      --  2 consecutive reads in case of write/read collision
        if (unsigned(axi_str_rxs_dpmem_rd_data_d1) = (rxs_mem_full_mask)) then
          rxs_axistream_next_state <= RESET_INIT_2; -- good to go fro second read
          AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_three_mask); --  rxs_mem_last_read_out_ptr rxs mem last
                                                          --  read out for write should be all 1's
        else
          rxs_axistream_next_state <= RESET_INIT_1; -- not init yet
          AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_three_mask); -- rxs_mem_last_read_out_ptr
        end if;

      when RESET_INIT_2 =>
      -- we must wait until the rx client interface has initialized the ptrs in dpmem
        if (unsigned(axi_str_rxs_dpmem_rd_data_d1) = (rxs_mem_full_mask)) then
          rxs_axistream_next_state <= READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_1; -- good to go
          AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_empty_mask); -- set address up for next state; read rxd_mem_next_available4write_ptr
        else
          rxs_axistream_next_state <= RESET_INIT_1; --  write/read collision may have occurred because we didn't
                                                    --  get same value twice
          AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_three_mask); -- rxs_mem_last_read_out_ptr
        end if;

      when READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_1 =>
        rxd_mem_next_available4write_ptr_1_cmb <= axi_str_rxs_dpmem_rd_data_d1(C_RXD_MEM_ADDR_WIDTH downto 0);
        rxs_axistream_next_state <= READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_2;
        AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_empty_mask); -- set address up for next state read; rxd_mem_next_available4write_ptr

      when READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_2 =>
        if (unsigned(axi_str_rxs_dpmem_rd_data_d1) = unsigned(rxd_mem_next_available4write_ptr_1_reg)) then -- good to go
          rxd_mem_next_available4write_ptr_cmb <= axi_str_rxs_dpmem_rd_data_d1(C_RXD_MEM_ADDR_WIDTH downto 0);
          rxs_axistream_next_state <= ADDR_SETUP_PAUSE_1;
          AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_two_mask); -- set address up for next state read;rxs_mem_next_available4write_ptr
        else
          AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_empty_mask); -- set address up for next state read; rxd_mem_next_available4write_ptr
          rxs_axistream_next_state <= READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_1; -- write/read collision may have occurred
                                                                               -- because we didn't get same value twice
        end if;

      when ADDR_SETUP_PAUSE_1 =>
        rxs_axistream_next_state <= READ_RXS_MEM_NEXT_AVAILABLE4WRITE_PTR_1;
        AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_two_mask); -- set address up for next state read;rxs_mem_next_available4write_ptr

      when READ_RXS_MEM_NEXT_AVAILABLE4WRITE_PTR_1 =>
        rxs_mem_next_available4write_ptr_1_cmb <= axi_str_rxs_dpmem_rd_data_d1(C_RXS_MEM_ADDR_WIDTH downto 0);
        rxs_axistream_next_state <= READ_RXS_MEM_NEXT_AVAILABLE4WRITE_PTR_2;
        AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_two_mask); -- set address up for next state read;rxs_mem_next_available4write_ptr

      when READ_RXS_MEM_NEXT_AVAILABLE4WRITE_PTR_2 =>
        if (unsigned(axi_str_rxs_dpmem_rd_data_d1) = unsigned(rxs_mem_next_available4write_ptr_1_reg)) then -- good to go
          rxs_mem_next_available4write_ptr_cmb <= axi_str_rxs_dpmem_rd_data_d1(C_RXS_MEM_ADDR_WIDTH downto 0);
          rxs_axistream_next_state <= ADDR_SETUP_PAUSE_2;
          AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_three_mask); -- set address up for next state read; rxs_mem_last_read_out_ptr
        else
          AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_two_mask); -- set address up for next state read;rxs_mem_next_available4write_ptr
          rxs_axistream_next_state <= READ_RXS_MEM_NEXT_AVAILABLE4WRITE_PTR_1;  --  write/read collision may have occurred
                                                                                --  because we didn't get same value twice
        end if;

      when ADDR_SETUP_PAUSE_2 =>
        rxs_axistream_next_state <= READ_RXS_MEM_LAST_READ_OUT_PTR;
        AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_three_mask); -- set address up for next state read; rxs_mem_last_read_out_ptr

      when READ_RXS_MEM_LAST_READ_OUT_PTR =>
      -- no need to double read this ptr, the other side does not write this location in memory
        if ((unsigned(axi_str_rxs_dpmem_rd_data_d1(C_RXS_MEM_ADDR_WIDTH downto 0)) = unsigned(rxs_mem_full_mask)) or (axi_str_rxs_dpmem_rd_data_d1(0) = 'X')) then -- to get rid of the xpm memory collision
          rxs_mem_last_read_out_ptr_cmb      <= rxs_mem_four_mask;
          rxs_mem_last_read_out_ptr_true_cmb <= std_logic_vector(rxs_mem_full_mask);
        else
          rxs_mem_last_read_out_ptr_cmb      <= unsigned(axi_str_rxs_dpmem_rd_data_d1(C_RXS_MEM_ADDR_WIDTH downto 0)) + 1;
          rxs_mem_last_read_out_ptr_true_cmb <= axi_str_rxs_dpmem_rd_data_d1(C_RXS_MEM_ADDR_WIDTH downto 0);
        end if;
        rxs_axistream_next_state  <= ADDR_SETUP_PAUSE_3;
        AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_one_mask); -- set address up for next state read; rxd_mem_last_read_out_ptr

      when ADDR_SETUP_PAUSE_3 =>
          rxs_axistream_next_state  <= READ_RXD_MEM_LAST_READ_OUT_PTR;
          AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_one_mask); -- set address up for next state read; rxd_mem_last_read_out_ptr

      when READ_RXD_MEM_LAST_READ_OUT_PTR =>
      -- no need to double read this ptr, the other side does not write this location in memory
        rxd_mem_last_read_out_ptr_cmb <= axi_str_rxs_dpmem_rd_data_d1(C_RXD_MEM_ADDR_WIDTH downto 0);
        if (rxs_mem_last_read_out_ptr_true_reg = std_logic_vector(rxs_mem_full_mask))then -- check to see if rxs mem is empty or ready to process
          if (rxs_mem_next_available4write_ptr_reg = std_logic_vector(rxs_mem_four_mask)) then -- rxs mem is empty
            rxs_axistream_next_state <= READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_1;
            AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_empty_mask); -- set address up for next state read; rxd_mem_next_available4write_ptr
          else -- rxs mem has a frame ready
            rxs_axistream_next_state <= PAUSE_READ_STATUS_WORD1;
            AXI_STR_RXS_DPMEM_ADDR   <= rxs_mem_last_read_out_ptr_reg; -- set address up for next state read; status word 1
          end if;
        else
          if (rxs_mem_next_available4write_ptr_reg = std_logic_vector(unsigned(rxs_mem_last_read_out_ptr_true_reg) + 1)) then -- rxs mem is empty
            rxs_axistream_next_state <= READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_1;
            AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_empty_mask); -- set address up for next state read; rxd_mem_next_available4write_ptr
          else -- rxs mem has a frame ready
            rxs_axistream_next_state <= PAUSE_READ_STATUS_WORD1;
            AXI_STR_RXS_DPMEM_ADDR   <= rxs_mem_last_read_out_ptr_reg; -- set address up for next state read; status word 1
          end if;
        end if;

      when PAUSE_READ_STATUS_WORD1 => -- delay so we can use register output of BRAM
         rxs_axistream_next_state <= READ_STATUS_WORD1;
         AXI_STR_RXS_DPMEM_ADDR   <= rxs_mem_last_read_out_ptr_reg; -- set address up for next state read; status word 1

      when READ_STATUS_WORD1 =>
        rxs_axistream_next_state  <= READ_STATUS_WORD2;
        rxs_mem_last_read_out_ptr_cmb <= rxs_mem_last_read_out_ptr_plus_one;
        rxs_mem_last_read_out_ptr_true_cmb <= rxs_mem_last_read_out_ptr_reg;
        AXI_STR_RXS_DPMEM_ADDR    <= std_logic_vector(rxs_mem_last_read_out_ptr_plus_one); -- set address up for next state read

      when READ_STATUS_WORD2 =>
        rxs_axistream_next_state  <= READ_STATUS_WORD3;
        rxs_mem_last_read_out_ptr_cmb <= rxs_mem_last_read_out_ptr_plus_one;
        rxs_mem_last_read_out_ptr_true_cmb <= rxs_mem_last_read_out_ptr_reg;
        AXI_STR_RXS_DPMEM_ADDR    <= std_logic_vector(rxs_mem_last_read_out_ptr_plus_one); -- set address up for next state read

      when READ_STATUS_WORD3 =>
        rxs_axistream_next_state  <= READ_STATUS_WORD4;
        rxs_mem_last_read_out_ptr_cmb <= rxs_mem_last_read_out_ptr_plus_one;
        rxs_mem_last_read_out_ptr_true_cmb <= rxs_mem_last_read_out_ptr_reg;
        AXI_STR_RXS_DPMEM_ADDR    <= std_logic_vector(rxs_mem_last_read_out_ptr_plus_one); -- set address up for next state read

      when READ_STATUS_WORD4 =>
        rxs_axistream_next_state  <= READ_STATUS_WORD5;
        rxs_mem_last_read_out_ptr_cmb <= rxs_mem_last_read_out_ptr_plus_one;
        rxs_mem_last_read_out_ptr_true_cmb <= rxs_mem_last_read_out_ptr_reg;
        AXI_STR_RXS_DPMEM_ADDR    <= std_logic_vector(rxs_mem_last_read_out_ptr_plus_one); -- set address up for next state read

      when READ_STATUS_WORD5 =>
        rxs_axistream_next_state  <= READ_STATUS_WORD6;
        rxs_mem_last_read_out_ptr_cmb <= rxs_mem_last_read_out_ptr_plus_one;
        rxs_mem_last_read_out_ptr_true_cmb <= rxs_mem_last_read_out_ptr_reg;
        AXI_STR_RXS_DPMEM_ADDR    <= std_logic_vector(rxs_mem_last_read_out_ptr_plus_one); -- set address up for next state read

      when READ_STATUS_WORD6 =>
        rxs_axistream_next_state  <= UPDATE_RXS_MEM_LAST_READ_OUT_PTR;
        AXI_STR_RXS_DPMEM_ADDR    <= std_logic_vector(rxs_mem_three_mask); -- set address up for next state read

      when UPDATE_RXS_MEM_LAST_READ_OUT_PTR =>
        rxs_axistream_next_state  <= SEND_STATUS_WORD1;
        AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_three_mask);
        AXI_STR_RXS_DPMEM_WR_DATA(35 downto C_RXS_MEM_ADDR_WIDTH + 1) <= (others => '0');
        AXI_STR_RXS_DPMEM_WR_DATA(C_RXS_MEM_ADDR_WIDTH downto 0) <= std_logic_vector(rxs_mem_last_read_out_ptr_cmb);
        AXI_STR_RXS_DPMEM_WR_EN(0)<= '1';
        rxs2rxd_frame_ready <= '1';

      when SEND_STATUS_WORD1 =>
        AXI_STR_RXS_VALID <= '1';
        AXI_STR_RXS_DATA  <= X"50000000";  --Set the flag,  all other bits are reserved
        rxs2rxd_frame_ready       <= '1';
        --  adding the following lines in case they process rxd before rxs and we end up stuck here,
        --  we update the pointers and memory
        if (rxd_addr_cntr_en = '1') then  --  update the read pointer for RXD memeory to free spaces up
                                          --  and as we send them over the RXD AXIStream
          rxd_mem_last_read_out_ptr_cmb <= std_logic_vector(rxd_mem_addr_cntr);
        end if;

        if (AXI_STR_RXS_READY = '1') then
          rxs_axistream_next_state  <= SEND_STATUS_WORD2;
        else
          rxs_axistream_next_state  <= SEND_STATUS_WORD1;
        end if;

      when SEND_STATUS_WORD2 =>
        AXI_STR_RXS_VALID <= '1';
        AXI_STR_RXS_DATA  <= rxs_status_word_2(31 downto 0);
        rxs2rxd_frame_ready       <= '1';

        --  adding the following lines in case they process rxd before rxs and we end up stuck here,
        --  we update the pointers and memory
        if (rxd_addr_cntr_en = '1') then  --  update the read pointer for RXD memeory to free spaces
                                          --  up and as we send them over the RXD AXIStream
          rxd_mem_last_read_out_ptr_cmb <= std_logic_vector(rxd_mem_addr_cntr);
        end if;

        if (AXI_STR_RXS_READY = '1') then
          rxs_axistream_next_state  <= SEND_STATUS_WORD3;
        else
          rxs_axistream_next_state  <= SEND_STATUS_WORD2;
        end if;

      when SEND_STATUS_WORD3 =>
        AXI_STR_RXS_VALID <= '1';
        AXI_STR_RXS_DATA  <= rxs_status_word_3(31 downto 0);
        rxs2rxd_frame_ready       <= '1';

        --  adding the following lines in case they process rxd before rxs and we end up stuck here,
        --  we update the pointers and memory
        if (rxd_addr_cntr_en = '1') then  --  update the read pointer for RXD memeory to free spaces
                                          --  up and as we send them over the RXD AXIStream
          rxd_mem_last_read_out_ptr_cmb <= std_logic_vector(rxd_mem_addr_cntr);
        end if;

        if (AXI_STR_RXS_READY = '1') then
          rxs_axistream_next_state  <= SEND_STATUS_WORD4;
        else
          rxs_axistream_next_state  <= SEND_STATUS_WORD3;
        end if;

      when SEND_STATUS_WORD4 =>
        AXI_STR_RXS_VALID <= '1';
        AXI_STR_RXS_DATA  <= rxs_status_word_4(31 downto 0);
        rxs2rxd_frame_ready       <= '1';

        --  adding the following  lines in case they process rxd before rxs and we end up stuck here,
        --  we update the pointers and memory
        if (rxd_addr_cntr_en = '1') then  --  update the read pointer for RXD memeory to free spaces up and
                                          --  as we send them over the RXD AXIStream
          rxd_mem_last_read_out_ptr_cmb <= std_logic_vector(rxd_mem_addr_cntr);
        end if;

        if (AXI_STR_RXS_READY = '1') then
          rxs_axistream_next_state  <= SEND_STATUS_WORD5;
        else
          rxs_axistream_next_state  <= SEND_STATUS_WORD4;
        end if;

      when SEND_STATUS_WORD5 =>
        AXI_STR_RXS_VALID <= '1';
        AXI_STR_RXS_DATA  <= rxs_status_word_5(31 downto 0);
        rxs2rxd_frame_ready       <= '1';

        --  adding the following lines in case they process rxd before rxs and we end up stuck here,
        --  we update the pointers and memory
        if (rxd_addr_cntr_en = '1') then  --  update the read pointer for RXD memeory to free spaces up and
                                          --  as we send them over the RXD AXIStream
          rxd_mem_last_read_out_ptr_cmb <= std_logic_vector(rxd_mem_addr_cntr);
        end if;

        if (AXI_STR_RXS_READY = '1') then
          rxs_axistream_next_state  <= SEND_STATUS_WORD6;
        else
          rxs_axistream_next_state  <= SEND_STATUS_WORD5;
        end if;

      when SEND_STATUS_WORD6 =>
        AXI_STR_RXS_VALID <= '1';
        AXI_STR_RXS_DATA  <= rxs_status_word_6(31 downto 0);
        AXI_STR_RXS_LAST  <= '1';
        rxs2rxd_frame_ready       <= '1';

        --  adding the following lines in case they process rxd before rxs and we end up stuck here,
        --  we update the pointers and memory
        if (rxd_addr_cntr_en = '1') then  --  update the read pointer for RXD memeory to free spaces up and
                                          --  as we send them over the RXD AXIStream
          rxd_mem_last_read_out_ptr_cmb <= std_logic_vector(rxd_mem_addr_cntr);
        end if;

        if (AXI_STR_RXS_READY = '1') then
          rxs_axistream_next_state  <= WAIT_FRAME_DONE;
        else
          rxs_axistream_next_state  <= SEND_STATUS_WORD6;
        end if;

      when WAIT_FRAME_DONE =>
        rxs2rxd_frame_ready <= '1';
        if (rxd_addr_cntr_en = '1') then  --  update the read pointer for RXD memeory to free spaces up and
                                          --  as we send them over the RXD AXIStream
          rxd_mem_last_read_out_ptr_cmb <= std_logic_vector(rxd_mem_addr_cntr);
        end if;
        if (rxd2rxs_frame_done = '0') then
          rxs_axistream_next_state  <= WAIT_FRAME_DONE;
        else
          rxs_axistream_next_state  <= UPDATE_RXD_MEM_LAST_READ_OUT_PTR;
        end if;

      when UPDATE_RXD_MEM_LAST_READ_OUT_PTR =>
        rxs_axistream_next_state <= REPEAT_AGAIN;

      when REPEAT_AGAIN =>
        rxs_axistream_next_state <= READ_RXD_MEM_NEXT_AVAILABLE4WRITE_PTR_1;
        AXI_STR_RXS_DPMEM_ADDR   <= std_logic_vector(rxs_mem_empty_mask); -- set address up for next state read

      when others   =>
        rxs_axistream_next_state         <= RESET_INIT_1;
    end case;
  end process;


    --------------------------------------------------------------------------
    -- receive data AXIStream State Machine
    -- RXDTSSM_REGS_PROCESS: registered process of the state machine
    -- RXDTSSM_CMB_PROCESS:  combinatorial next-state logic
    -- ETHIP-4375: Added 2 Extra states to state machine:
    --  1.WRITE_FIRST_WORD -> Write the first word to FIFO
    -- 	2.LOAD_FIRST_WORD  -> Load First word to fifoDataOut_1d
    -- ETHIP-4543: Added Extra condition to deassert fifo_wr_en as soon as all
    -- the words of the frame are written to fifo and exit RD_FRAME_FROM_MEM state
    -- if (rxd_word_cnt = frame_length_words)
    --------------------------------------------------------------------------

    RXDTSSM_REGS_PROCESS: process (AXI_STR_RXD_ACLK)
    begin
      if rising_edge(AXI_STR_RXD_ACLK) then
        if(RESET2AXI_STR_RXD='1' or RESET2AXI_STR_RXS='1') then
          rxd_axistream_current_state <= IDLE;
        else
          rxd_axistream_current_state <= rxd_axistream_next_state;
        end if;
      end if;
    end process;

    fifoEmpty_1d_PROCESS: process (AXI_STR_RXD_ACLK)
    begin
      if rising_edge(AXI_STR_RXD_ACLK) then
          fifoEmpty_1d <= fifoEmpty;
      end if;
    end process;

    fifoDataOut_1d_PROCESS: process (AXI_STR_RXD_ACLK)
    begin
      if rising_edge(AXI_STR_RXD_ACLK) then
          if (fifoRdEn = '1') then
             fifoDataOut_1d <= fifoDataOut;
          end if;
      end if;
    end process;

    LAST_READY_LATCH_PROCESS : process (AXI_STR_RXD_ACLK)
    begin
      if rising_edge(AXI_STR_RXD_ACLK) then
         AXI_STR_RXD_READY_1D <= AXI_STR_RXD_READY;
         if (AXI_STR_RXD_READY_RED = '1') then
            LAST_READY_DEASSERT_LATCH <= '0';
         elsif (LAST_READY_DEASSERT = '1') then
            LAST_READY_DEASSERT_LATCH <= '1';
         end if;
      end if;
    end process;
    AXI_STR_RXD_READY_RED <= AXI_STR_RXD_READY and (not(AXI_STR_RXD_READY_1D));
    LAST_READY_DEASSERT   <= AXI_STR_RXD_LAST_INT and (not(AXI_STR_RXD_READY));

    AXI_STR_LAST_1D_PROCESS : process (AXI_STR_RXD_ACLK)
    begin
      if rising_edge(AXI_STR_RXD_ACLK) then
         AXI_STR_RXD_LAST_INT_1D <= AXI_STR_RXD_LAST_INT;
      end if;
    end process;
    AXI_STR_RXD_LAST_FED <= (not(AXI_STR_RXD_LAST_INT)) and AXI_STR_RXD_LAST_INT_1D;

    AXI_STR_LAST_LATCH : process (AXI_STR_RXD_ACLK)
    begin
      if rising_edge(AXI_STR_RXD_ACLK) then
         if (fifoEmpty = '0') then
            AXI_STR_RXD_LAST_FALL_LATCH <= '0';
         elsif (AXI_STR_RXD_LAST_FED = '1') then
            AXI_STR_RXD_LAST_FALL_LATCH <= '1';
         end if;
      end if;
    end process;

    AXI_STR_STRB_CHK_GEN : process (AXI_STR_RXD_ACLK)
    begin
      if rising_edge(AXI_STR_RXD_ACLK) then
         if (fifoRdEn = '1') then
            AXI_STR_RXD_STRB_CHK <= '0';
         elsif (AXI_STR_RXD_LAST_FALL_LATCH = '1') then
            AXI_STR_RXD_STRB_CHK <= '1';
         elsif (AXI_STR_RXD_READY_RED = '1') then
            AXI_STR_RXD_STRB_CHK <= '0';
         end if;
      end if;
    end process;

    RXDTSSM_CMB_PROCESS: process (
      rxd_axistream_current_state,
      rxs2rxd_frame_ready,
      AXI_STR_RXD_READY,
      frame_length_words,
      rxd_word_cnt,
      rxd_addr_cntr_load,
      fifoEmpty,
      fifoEmpty_1d,
      fifoAlmostFull,
      AXI_STR_RXD_LAST_FALL_LATCH,
      rxd2rxs_frame_done,
      rxs2rxd_frame_done
      )
    begin

    case rxd_axistream_current_state is

      when IDLE =>
        if(rxs2rxd_frame_ready = '1' and rxd2rxs_frame_done = '0') then
          rxd_axistream_next_state <= PRIME;
        else
          rxd_axistream_next_state <= IDLE;
        end if;

      when PRIME =>
        rxd_axistream_next_state <= WRITE_FIRST_WORD;
        
      when WRITE_FIRST_WORD =>
	rxd_axistream_next_state <= LOAD_FIRST_WORD;
	
      when LOAD_FIRST_WORD =>
	if (fifoEmpty = '0') then
	  rxd_axistream_next_state <= RD_FRAME_FROM_MEM;
	else
	  rxd_axistream_next_state <= LOAD_FIRST_WORD;
	end if;  
	
      when RD_FRAME_FROM_MEM =>
        if (((rxd_word_cnt = frame_length_words - 1) or (rxd_word_cnt = frame_length_words)) and fifoEmpty_1d = '0') then -- ETHIP-4543
          rxd_axistream_next_state <= WAIT_END_FRAME;
        elsif (fifoAlmostFull = '1') then
          rxd_axistream_next_state <= ALMOST_FULL_WAIT1;
        else
          rxd_axistream_next_state <= RD_FRAME_FROM_MEM;
        end if;

      when ALMOST_FULL_WAIT1 =>
        rxd_axistream_next_state <= ALMOST_FULL_WAIT2;

      when ALMOST_FULL_WAIT2 =>
        if (fifoAlmostFull = '0') then
          rxd_axistream_next_state <= ALMOST_FULL_WAIT3;
        else
          rxd_axistream_next_state <= ALMOST_FULL_WAIT2;
        end if;

      when ALMOST_FULL_WAIT3 =>
        rxd_axistream_next_state <= ALMOST_FULL_WAIT4;

      when ALMOST_FULL_WAIT4 =>
        rxd_axistream_next_state <= RD_FRAME_FROM_MEM;

      when WAIT_END_FRAME =>
        if (AXI_STR_RXD_LAST_FALL_LATCH = '1') then
          rxd_axistream_next_state <= PRE_IDLE;
        else
          rxd_axistream_next_state <= WAIT_END_FRAME;
        end if;

      when PRE_IDLE =>
        if (rxs2rxd_frame_done = '0') then
          rxd_axistream_next_state  <= PRE_IDLE;
        else
          rxd_axistream_next_state  <= IDLE;
        end if;

      when others   =>
        rxd_axistream_next_state <= IDLE;

    end case;
  end process;

  rxd_addr_cntr_en    <= '1' when ((fifoWrEn = '1') and (fifoAlmostFull = '0') and
                                   (rxd_word_cnt < frame_length_words - 1)) else
                         '1' when ((rxd_axistream_current_state = ALMOST_FULL_WAIT4) and (fifoAlmostFull = '0') and
                                   (rxd_word_cnt < frame_length_words - 1)) else
                         '1' when ((rxd_axistream_current_state = PRIME)) else
                         '0';

  AXI_STR_RXD_DPMEM_ADDR <= std_logic_vector(rxd_mem_addr_cntr);

  fifoWrEn            <= '1' when ((rxd_axistream_current_state = RD_FRAME_FROM_MEM) and
                                   (rxd_word_cnt < frame_length_words)) else     -- ETHIP-4543         
                         '1' when (rxd_axistream_current_state = WRITE_FIRST_WORD) else
                         '1' when ((rxd_axistream_current_state = LOAD_FIRST_WORD) and 
                                   (rxd_word_cnt < frame_length_words)) else
                         '0';

  fifoDataIn          <= AXI_STR_RXD_DPMEM_RD_DATA(35 downto 0);

  rxd2rxs_frame_done  <= '1' when (rxd_axistream_current_state = PRE_IDLE) else
                         '0';

  rxs2rxd_frame_done  <= '1' when (rxs_axistream_current_state = WAIT_FRAME_DONE) else
                         '0';

  rxd_addr_cntr_load  <= '1' when (rxd_axistream_current_state = IDLE) else
                         '0';

  fifoRdEn            <= '1' when ((rxd_axistream_current_state = LOAD_FIRST_WORD and fifoEmpty = '0') or (AXI_STR_RXD_READY = '1')  or (RESET2AXI_STR_RXD = '1')) else
                         '0';
  AXI_STR_RXD_DATA    <= fifoDataOut_1d(4 to 35);
  AXI_STR_RXD_VALID   <=  '1' when (LAST_READY_DEASSERT_LATCH = '1') else 
                          not(fifoEmpty_1d);
  AXI_STR_RXD_STRB    <= "0000" when (AXI_STR_RXD_STRB_CHK = '1') else
                         fifoDataOut_1d(0 to 3);
  AXI_STR_RXD_LAST_INT <= '1' when ((rxd_axistream_current_state = WAIT_END_FRAME and fifoEmpty = '1' and fifoDataCount = "000001") or (LAST_READY_DEASSERT_LATCH = '1')) else
                          '0';
  AXI_STR_RXD_LAST     <= AXI_STR_RXD_LAST_INT;

  COUNT_RXD_WORDS_READ : process (AXI_STR_RXD_ACLK)
  begin
    if rising_edge(AXI_STR_RXD_ACLK) then
      if RESET2AXI_STR_RXD = '1' then
        rxd_word_cnt   <= 0;
      else
        if (rxd_axistream_current_state = IDLE or rxd_word_cnt = 32767) then
          rxd_word_cnt   <= 0;
        elsif (fifoWrEn = '1') then
          rxd_word_cnt <= rxd_word_cnt + 1;
        end if;
      end if;
    end if;
  end process;

  DETECT_FIFO_ALMOST_FULL : process(fifoDataCount, fifoEmpty_1d)
  begin
    fifoAlmostFull  <= '0';
    if(to_integer(unsigned(fifoDataCount))>28 and fifoEmpty_1d='0') then
      fifoAlmostFull <= '1';
    end if;
  end process;


----  Since this fifo is removed during proc_common re-factoring. Taking this module into buffer.
---------------------------------------------------------------------
  --- removing this fifo as it is lo longer supported by the proc common . Using lib_fifo instead which is recommended.
  ELASTIC_FIFO : basic_sfifo_fg
  generic map(
    C_DWIDTH                      => 36,
      -- FIFO data Width (Read and write data ports are symetric)
    C_DEPTH                       => 32,
      -- FIFO Depth (set to power of 2)
    C_HAS_DATA_COUNT              => 1,
      -- 0 = DataCount not used
      -- 1 = Data Count used
    C_DATA_COUNT_WIDTH            => 6,
    -- Data Count bit width (Max value is log2(C_DEPTH))
    C_IMPLEMENTATION_TYPE         => 0,
      --  0 = Common Clock BRAM / Distributed RAM (Synchronous FIFO)
      --  1 = Common Clock Shift Register (Synchronous FIFO)
    C_MEMORY_TYPE                 => 2,
      --   0 = Any
      --   1 = BRAM
      --   2 = Distributed Memory
      --   3 = Shift Registers
    C_PRELOAD_REGS                => 1,
      -- 0 = normal
      -- 1 for FWFT
    C_PRELOAD_LATENCY             => 0,
      -- 0 for FWFT
      -- 1 = normal
    C_USE_FWFT_DATA_COUNT         => 1,
      -- 0 = normal
      -- 1 for FWFT
    C_FAMILY                      =>  C_FAMILY
    )
  port map(
    CLK                           =>  AXI_STR_RXD_ACLK,
    DIN                           =>  fifoDataIn,
    RD_EN                         =>  fifoRdEn,
    SRST                          =>  RESET2AXI_STR_RXD,
    WR_EN                         =>  fifoWrEn,
    DATA_COUNT                    =>  fifoDataCount,
    DOUT                          =>  fifoDataOut,
    EMPTY                         =>  fifoEmpty,
    FULL                          =>  fifoFull
    );

---  ELASTIC_FIFO : entity lib_fifo_v1_0.sync_fifo_fg
---  generic map(
---    C_DCOUNT_WIDTH     => 6,
---    C_HAS_DCOUNT       => 1,
---    C_MEMORY_TYPE      => 0,
---    C_PRELOAD_LATENCY  => 0,
---    C_PRELOAD_REGS     => 1,
---    C_READ_DATA_WIDTH  => 36,
---    C_READ_DEPTH       => 32,
---    C_WRITE_DATA_WIDTH => 36,
---    C_WRITE_DEPTH      => 32,
---    C_FAMILY           => C_FAMILY
---    )
---  port map(
---    Clk         => AXI_STR_RXD_ACLK,----- : in  std_logic;
---    Sinit       => RESET2AXI_STR_RXD,----- : in  std_logic;
---    Din         => fifoDataIn,----- : in  std_logic_vector(C_WRITE_DATA_WIDTH-1 downto 0);
---    Wr_en       => fifoWrEn,----- : in  std_logic;
---    Rd_en       => fifoRdEn,----- : in  std_logic;
---    Dout        => fifoDataOut,----- : out std_logic_vector(C_READ_DATA_WIDTH-1 downto 0);
---    Almost_full => OPEN,----- : out std_logic;
---    Full        => fifoFull,----- : out std_logic;
---    Empty       => fifoEmpty,----- : out std_logic;
---    Rd_ack      => OPEN,----- : out std_logic;
---    Wr_ack      => OPEN,----- : out std_logic;
---    Rd_err      => OPEN,----- : out std_logic;
---    Wr_err      => OPEN,----- : out std_logic;
---    Data_count  => fifoDataCount ----- : out std_logic_vector(C_DCOUNT_WIDTH-1 downto 0)
---    );

end rtl;


------------------------------------------------------------------------
-- Title      : Package for the registers_pack logic
-- Project    : Tri-Mode Ethernet FIFO
------------------------------------------------------------------------
-- File       : registers_pack.vhd
-- Author     : Xilinx Inc.
------------------------------------------------------------------------
-- (c) Copyright 2012 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
------------------------------------------------------------------------
-- Description:  This package contains all component declarations for
--               the entiries which make up the Register logic
------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;



package registers_pack is

  component registers
  generic
  (
    C_FAMILY       : string   := "virtex5";
    C_TXVLAN_TRAN  : integer  := 1;
    C_TXVLAN_TAG   : integer  := 1;
    C_TXVLAN_STRP  : integer  := 1;
    C_RXVLAN_TRAN  : integer  := 1;
    C_RXVLAN_TAG   : integer  := 1;
    C_RXVLAN_STRP  : integer  := 1;
    C_MCAST_EXTEND : integer  := 1;
    C_TXVLAN_WIDTH : integer  := 1;
    C_RXVLAN_WIDTH : integer  := 1
  );
  port
  (
    AxiClk                    : in  std_logic;                    --  AXI4-Lite Clock
    AXI_STR_TXD_ACLK          : in  std_logic;                    --  AXI-Stream Transmit Data Clock
    RxClClk                   : in  std_logic;                    --  Receive Client Clock
    AxiReset                  : in  std_logic;                    --  AXI4-Lite Reset
    IP2Bus_Data               : out std_logic_vector(0 to 31);    --  AXI Ethernet to AXI4-Lite Data
    IP2Bus_WrAck              : out std_logic;                    --  AXI Ethernet to AXI4-Lite Write Ack
    IP2Bus_RdAck              : out std_logic;                    --  AXI Ethernet to AXI4-Lite Read Ack
    Bus2IP_Addr               : in  std_logic_vector(0 to 31);    --  AXI4-Lite to AXI Ethernet Addr
    Bus2IP_Data               : in  std_logic_vector(0 to 31);    --  AXI4-Lite to AXI Ethernet Data
    Bus2IP_RNW                : in  std_logic;                    --  AXI4-Lite to AXI Ethernet RNW
    Bus2IP_CS                 : in  std_logic_vector(0 to 10);    --  AXI4-Lite to AXI Ethernet CS
    Bus2IP_RdCE               : in  std_logic_vector(0 to 41);    --  AXI4-Lite to AXI Ethernet RdCE
    Bus2IP_WrCE               : in  std_logic_vector(0 to 41);    --  AXI4-Lite to AXI Ethernet WrCE
    IntrptsIn                 : in  std_logic_vector(23 to 31);   --  Interrupts in
    TPReq                     : out std_logic;                    --  Transmit Pause Request
    CrRegData                 : out std_logic_vector(17 to 31);   --  RAF Register
    TpRegData                 : out std_logic_vector(16 to 31);   --  Transmit Pause Data
    IfgpRegData               : out std_logic_vector(24 to 31);   --  Inter Frame Gap Data
    IsRegData                 : out std_logic_vector(23 to 31);   --  Interrupt Status Register
    IpRegData                 : out std_logic_vector(23 to 31);   --  Interrupt Pending Register
    IeRegData                 : out std_logic_vector(23 to 31);   --  Interrupt Enable Register
    IntrptOut                 : out std_logic;                    --  Interrupt Out
    TtagRegData               : out std_logic_vector(0 to 31);    --  Transmit Tag Register
    RtagRegData               : out std_logic_vector(0 to 31);    --  Receive Tag Register
    Tpid0RegData              : out std_logic_vector(0 to 31);    --  VLAN TPID Reg 0
    Tpid1RegData              : out std_logic_vector(0 to 31);    --  VLAN TPID Reg 1
    pcspma_status_cross       : in  std_logic_vector(16 to 31);   --  PCS PMA Link Status Vector
    UawLRegData               : out std_logic_vector(0 to 31);    --  Unicast Address Word Lower
    UawURegData               : out std_logic_vector(16 to 31);   --  Unicast Address Word Upper
    RxClClkMcastAddr          : in  std_logic_vector(0 to 14);    --  Receive Extended Multicast Address
    RxClClkMcastEn            : in  std_logic;                    --  Receive Extended Multicast Enable
    RxClClkMcastRdData        : out std_logic_vector(0 to 0);     --  Receive Extended Multicast Data
    AxiStrTxDClkTxVlanAddr    : in  std_logic_vector(0 to 11);    --  Transmit VLAN BRAM Addr
    AxiStrTxDClkTxVlanRdData  : out std_logic_vector(18 to 31);   --  Transmit VLAN BRAM Read Data
    RxClClkRxVlanAddr         : in  std_logic_vector(0 to 11);    --  Receive VLAN BRAM Addr
    RxClClkRXVlanRdData       : out std_logic_vector(18 to 31);   --  Receive VLAN BRAM Read Data
    AxiStrTxDClkTxVlanBramEnA : in  std_logic;                    --  Transmit VLAN BRAM Enable
    RxClClkRxVlanBramEnA      : in  std_logic                     --  Receive VLAN BRAM Enable
  );
  end component;


  component reg_tp
    port    (
             Clk      : in  std_logic;                  --  Clk     in
             RST      : in  std_logic;                  --  RST     in
             RdCE     : in  std_logic;                  --  RdCE    in
             WrCE     : in  std_logic;                  --  WrCE    in
             DataIn   : in  std_logic_vector(16 to 31); --  DataIn  in
             DataOut  : out std_logic_vector(16 to 31); --  DataOut out
             RegData  : out std_logic_vector(16 to 31); --  RegData out
             TPReq    : out std_logic                   --  TPReq   out
            );
  end component;


  component reg_is
    port    (
             Clk      : in  std_logic;                      --Clk      in
             RST      : in  std_logic;                      --RST      in
             RdCE     : in  std_logic;                      --RdCE     in
             WrCE     : in  std_logic;                      --WrCE     in
             Intrpts  : in  std_logic_vector(23 to 31);     --Intrpts  in
             DataIn   : in  std_logic_vector(23 to 31);     --DataIn   in
             DataOut  : out std_logic_vector(23 to 31);     --DataOut  out
             RegData  : out std_logic_vector(23 to 31)      --RegData  out
            );
  end component;


  component reg_ip
    port    (
             Clk      : in  std_logic;                    --  Clk Input
             RST      : in  std_logic;                    --  RST Input
             RdCE     : in  std_logic;                    --  RdCE Input
             IsIn     : in std_logic_vector(23 to 31);    --  IsIn Input
             IeIn     : in std_logic_vector(23 to 31);    --  IeIn Input
             DataOut  : out std_logic_vector(23 to 31);   --  DataOut Output
             RegData  : out std_logic_vector(23 to 31);   --  RegData Output
             Intrpt   : out std_logic                     --  Intrpt Output
            );
  end component;


  component reg_16bl
    port    (
             Clk      : in  std_logic;                      --  Clk Input
             RST      : in  std_logic;                      --  RST Input
             RdCE     : in  std_logic;                      --  RdCE Input
             WrCE     : in  std_logic;                      --  WrCE Input
             DataIn   : in  std_logic_vector(16 to 31);     --  DataIn Input
             DataOut  : out std_logic_vector(16 to 31);     --  DataOut Output
             RegData  : out std_logic_vector(16 to 31);     --  RegData Output
             TPReq    : out std_logic                       --  TPReq Output
            );
  end component;


  component reg_32b
    port    (
             Clk      : in  std_logic;                      --  Clk Input
             RST      : in  std_logic;                      --  RST Input
             RdCE     : in  std_logic;                      --  RdCE Input
             WrCE     : in  std_logic;                      --  WrCE Input
             DataIn   : in  std_logic_vector(0 to 31);      --  DataIn Input
             DataOut  : out std_logic_vector(0 to 31);      --  DataOut Output
             RegData  : out std_logic_vector(0 to 31);      --  RegData Output
             TPReq    : out std_logic                       --  TPReq Output
            );
  end component;


  component reg_cr
    port    (
             Clk      : in  std_logic;  --intPlbClk               --  Clk        in
                                                                  --
             RST      : in  std_logic;                            --  RST        in
             RdCE     : in  std_logic;                            --  RdCE       in
             WrCE     : in  std_logic;                            --  WrCE       in
             DataIn   : in  std_logic_vector(17 to 31);           --  DataIn     in
             DataOut  : out std_logic_vector(17 to 31);           --  DataOut    out
             RegData  : out std_logic_vector(17 to 31)            --  RegData    out
            );
  end component;


  component reg_ie
    port    (
             Clk      : in  std_logic;                    --  Clk Input
             RST      : in  std_logic;                    --  RST Input
             RdCE     : in  std_logic;                    --  RdCE Input
             WrCE     : in  std_logic;                    --  WrCE Input
             DataIn   : in  std_logic_vector(23 to 31);   --  DataIn Input
             DataOut  : out std_logic_vector(23 to 31);   --  DataOut Output
             RegData  : out std_logic_vector(23 to 31)    --  RegData Output
            );
  end component;


  component reg_ifgp
    port    (
             Clk      : in  std_logic;                  --  Clk Input
             RST      : in  std_logic;                  --  RST Input
             RdCE     : in  std_logic;                  --  RdCE Input
             WrCE     : in  std_logic;                  --  WrCE Input
             DataIn   : in  std_logic_vector(24 to 31); --  DataIn Input
             DataOut  : out std_logic_vector(24 to 31); --  DataOut Output
             RegData  : out std_logic_vector(24 to 31)  --  RegData Output
            );
  end component;


end registers_pack;


------------------------------------------------------------------------------
-- $Id: reg_tp.vhd,v 1.1.2.2 2010/12/15 22:53:05 mwelter Exp $
------------------------------------------------------------------------------
-- reg_tp - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        reg_tp.vhd
-- Version:         v1.01a
-- Description:     Include a meaningful description of your file. Multi-line
--                  descriptions should align with each other
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:
-- History:
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.registers_pack.all;

entity reg_tp is
    port    (
             Clk      : in  std_logic;                  --  Clk     in
             RST      : in  std_logic;                  --  RST     in
             RdCE     : in  std_logic;                  --  RdCE    in
             WrCE     : in  std_logic;                  --  WrCE    in
             DataIn   : in  std_logic_vector(16 to 31); --  DataIn  in
             DataOut  : out std_logic_vector(16 to 31); --  DataOut out
             RegData  : out std_logic_vector(16 to 31); --  RegData out
             TPReq    : out std_logic                   --  TPReq   out
            );
end reg_tp;

------------------------------------------------------------------------------
-- Architecture
------------------------------------------------------------------------------

architecture imp of reg_tp is

------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

signal reg_data : std_logic_vector(16 to 31);
signal wrCE_d   : std_logic;

begin

------------------------------------------------------------------------------
-- Concurrent Signal Assignments
------------------------------------------------------------------------------

RegData   <= reg_data;

------------------------------------------------------------------------------
-- BUS_READ_PROCESS
------------------------------------------------------------------------------

BUS_READ_PROCESS : process (RdCE, reg_data)
begin
    for i in 16 to 31
    loop
        DataOut(i) <= RdCE and reg_data(i);
    end loop;
end process;

------------------------------------------------------------------------------
-- BUS_WRITE_PROCESS
------------------------------------------------------------------------------

BUS_WRITE_PROCESS : process (Clk)
begin
    if (Clk'event and Clk = '1')
    then
        if (Rst = '1') then
          reg_data <= (others => '0');
          TPReq    <= '0';
          wrCE_d   <= '0';
        elsif (WrCE = '1') then
          reg_data <= DataIn;
          TPReq    <= wrCE_d;
          wrCE_d   <= WrCE;
        else
          TPReq    <= wrCE_d;
          wrCE_d   <= WrCE;
        end if;
    end if;
end process;

end imp;


------------------------------------------------------------------------------
-- reg_is - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        reg_is.vhd
-- Version:         v1.01a
-- Description:     Include a meaningful description of your file. Multi-line
--                  descriptions should align with each other
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:
-- History:
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.registers_pack.all;

entity reg_is is
    port    (
             Clk      : in  std_logic;                      --Clk      in
             RST      : in  std_logic;                      --RST      in
             RdCE     : in  std_logic;                      --RdCE     in
             WrCE     : in  std_logic;                      --WrCE     in
             Intrpts  : in  std_logic_vector(23 to 31);     --Intrpts  in
             DataIn   : in  std_logic_vector(23 to 31);     --DataIn   in
             DataOut  : out std_logic_vector(23 to 31);     --DataOut  out
             RegData  : out std_logic_vector(23 to 31)      --RegData  out
            );
end reg_is;

------------------------------------------------------------------------------
-- Architecture
------------------------------------------------------------------------------

architecture imp of reg_is is

------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

signal reg_data : std_logic_vector(23 to 31);

begin

------------------------------------------------------------------------------
-- Concurrent Signal Assignments
------------------------------------------------------------------------------

RegData   <= reg_data;

------------------------------------------------------------------------------
-- BUS_READ_PROCESS
------------------------------------------------------------------------------

BUS_READ_PROCESS : process (RdCE, reg_data)
begin
    for i in 23 to 31 loop
        DataOut(i) <= RdCE and reg_data(i);
    end loop;
end process;

------------------------------------------------------------------------------
-- BUS_WRITE_PROCESS
------------------------------------------------------------------------------

BUS_WRITE_PROCESS : process (Clk)
begin
    if (Clk'event and Clk = '1') then
      for i in 23 to 31 loop
        if (Rst = '1') then
          reg_data(i) <= '0';
        elsif (WrCE = '1' and DataIn(i) = '1') then
          reg_data(i) <= '0';
        elsif (Intrpts(i) = '1') then
          reg_data(i) <= '1';
        else
          null;
        end if;
      end loop;
    end if;
end process;

end imp;


------------------------------------------------------------------------------
-- reg_ip - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        reg_ip.vhd
-- Version:         v1.01a
-- Description:     Include a meaningful description of your file. Multi-line
--                  descriptions should align with each other
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:
-- History:
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.registers_pack.all;

entity reg_ip is
    port    (
             Clk      : in  std_logic;                    --  Clk Input
             RST      : in  std_logic;                    --  RST Input
             RdCE     : in  std_logic;                    --  RdCE Input
             IsIn     : in std_logic_vector(23 to 31);    --  IsIn Input
             IeIn     : in std_logic_vector(23 to 31);    --  IeIn Input
             DataOut  : out std_logic_vector(23 to 31);   --  DataOut Output
             RegData  : out std_logic_vector(23 to 31);   --  RegData Output
             Intrpt   : out std_logic                     --  Intrpt Output
            );
end reg_ip;

------------------------------------------------------------------------------
-- Architecture
------------------------------------------------------------------------------

architecture imp of reg_ip is

------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

signal reg_data : std_logic_vector(23 to 31);

begin

------------------------------------------------------------------------------
-- Concurrent Signal Assignments
------------------------------------------------------------------------------

RegData   <= reg_data;

------------------------------------------------------------------------------
-- BUS_READ_PROCESS
------------------------------------------------------------------------------

BUS_READ_PROCESS : process (RdCE, reg_data)
begin
    for i in 23 to 31
    loop
        DataOut(i) <= RdCE and reg_data(i);
    end loop;
end process;

BUS_WRITE_PROCESS : process (Clk, IsIn, IeIn)
begin
  if (Clk'event and Clk = '1') then
    if (Rst = '1') then
      reg_data <= (others => '0');
      Intrpt   <= '0';
    else
      reg_data <= IsIn and IeIn;
      if (reg_data = "000000000") then
        Intrpt   <= '0';
      else
        Intrpt   <= '1';
      end if;
    end if;
  end if;
end process;

end imp;


------------------------------------------------------------------------------
-- $Id: reg_ifgp.vhd,v 1.1.2.2 2010/12/15 22:53:05 mwelter Exp $
------------------------------------------------------------------------------
-- reg_ifgp - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        reg_ifgp.vhd
-- Version:         v1.01a
-- Description:     Include a meaningful description of your file. Multi-line
--                  descriptions should align with each other
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:
-- History:
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.registers_pack.all;

entity reg_ifgp is
    port    (
             Clk      : in  std_logic;                  --  Clk Input
             RST      : in  std_logic;                  --  RST Input
             RdCE     : in  std_logic;                  --  RdCE Input
             WrCE     : in  std_logic;                  --  WrCE Input
             DataIn   : in  std_logic_vector(24 to 31); --  DataIn Input
             DataOut  : out std_logic_vector(24 to 31); --  DataOut Output
             RegData  : out std_logic_vector(24 to 31)  --  RegData Output
            );
end reg_ifgp;

------------------------------------------------------------------------------
-- Architecture
------------------------------------------------------------------------------

architecture imp of reg_ifgp is

------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

signal reg_data : std_logic_vector(24 to 31);

begin

------------------------------------------------------------------------------
-- Concurrent Signal Assignments
------------------------------------------------------------------------------

RegData   <= reg_data;

------------------------------------------------------------------------------
-- BUS_READ_PROCESS
------------------------------------------------------------------------------

BUS_READ_PROCESS : process (RdCE, reg_data)
begin
    for i in 24 to 31
    loop
        DataOut(i) <= RdCE and reg_data(i);
    end loop;
end process;

------------------------------------------------------------------------------
-- BUS_WRITE_PROCESS
------------------------------------------------------------------------------

BUS_WRITE_PROCESS : process (Clk)
begin
    if (Clk'event and Clk = '1')
    then
        if (Rst = '1')
        then
            reg_data <= (others => '0');
        elsif (WrCE = '1')
        then
            reg_data <= DataIn;
        end if;
    end if;
end process;

end imp;


------------------------------------------------------------------------------
-- reg_ie - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        reg_ie.vhd
-- Version:         v1.01a
-- Description:     Include a meaningful description of your file. Multi-line
--                  descriptions should align with each other
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:
-- History:
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.registers_pack.all;

entity reg_ie is
    port    (
             Clk      : in  std_logic;                    --  Clk Input
             RST      : in  std_logic;                    --  RST Input
             RdCE     : in  std_logic;                    --  RdCE Input
             WrCE     : in  std_logic;                    --  WrCE Input
             DataIn   : in  std_logic_vector(23 to 31);   --  DataIn Input
             DataOut  : out std_logic_vector(23 to 31);   --  DataOut Output
             RegData  : out std_logic_vector(23 to 31)    --  RegData Output
            );
end reg_ie;

------------------------------------------------------------------------------
-- Architecture
------------------------------------------------------------------------------

architecture imp of reg_ie is

------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

signal reg_data : std_logic_vector(23 to 31);

begin

------------------------------------------------------------------------------
-- Concurrent Signal Assignments
------------------------------------------------------------------------------

RegData   <= reg_data;

------------------------------------------------------------------------------
-- BUS_READ_PROCESS
------------------------------------------------------------------------------

BUS_READ_PROCESS : process (RdCE, reg_data)
begin
    for i in 23 to 31
    loop
        DataOut(i) <= RdCE and reg_data(i);
    end loop;
end process;

------------------------------------------------------------------------------
-- BUS_WRITE_PROCESS
------------------------------------------------------------------------------

BUS_WRITE_PROCESS : process (Clk)
begin
    if (Clk'event and Clk = '1')
    then
        if (Rst = '1')
        then
            reg_data <= (others => '0');
        elsif (WrCE = '1')
        then
            reg_data <= DataIn;
        end if;
    end if;
end process;

end imp;


------------------------------------------------------------------------------
-- reg_cr - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        reg_cr.vhd
-- Version:         v1.01a
-- Description:     Include a meaningful description of your file. Multi-line
--                  descriptions should align with each other
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:
-- History:
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.registers_pack.all;

entity reg_cr is
    port    (
             Clk      : in  std_logic;  --intPlbClk               --  Clk        in
                                                                  --
             RST      : in  std_logic;                            --  RST        in
             RdCE     : in  std_logic;                            --  RdCE       in
             WrCE     : in  std_logic;                            --  WrCE       in
             DataIn   : in  std_logic_vector(17 to 31);           --  DataIn     in
             DataOut  : out std_logic_vector(17 to 31);           --  DataOut    out
             RegData  : out std_logic_vector(17 to 31)            --  RegData    out
            );
end reg_cr;

------------------------------------------------------------------------------
-- Architecture
------------------------------------------------------------------------------

architecture imp of reg_cr is

------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

signal reg_data : std_logic_vector(17 to 31);

begin

------------------------------------------------------------------------------
-- Concurrent Signal Assignments
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- REG_DATA_PROCESS
------------------------------------------------------------------------------

REG_DATA_PROCESS : process (reg_data)
begin
  for i in 17 to 31 loop
      RegData(i) <= reg_data(i);
  end loop;
end process;

------------------------------------------------------------------------------
-- BUS_READ_PROCESS
------------------------------------------------------------------------------

BUS_READ_PROCESS : process (RdCE, reg_data)
begin
  for i in 17 to 31 loop
     DataOut(i) <= RdCE and reg_data(i);
  end loop;
end process;

------------------------------------------------------------------------------
-- BUS_WRITE_PROCESS
------------------------------------------------------------------------------

BUS_WRITE_PROCESS : process (Clk)
begin
    if (Clk'event and Clk = '1')
    then
        if (Rst = '1')
        then
            reg_data <= (others => '0');
        elsif (WrCE = '1')
        then
            reg_data(17)       <= DataIn(17);
            reg_data(19 to 30) <= DataIn(19 to 30);
            reg_data(18)       <= '0';
            reg_data(31)       <= '0';
        end if;
    end if;
end process;

end imp;


------------------------------------------------------------------------------
-- $Id: reg_32b.vhd,v 1.1.2.2 2010/12/15 22:53:05 mwelter Exp $
------------------------------------------------------------------------------
-- reg_32b - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        reg_32b.vhd
-- Version:         v2.00a
-- Description:     Include a meaningful description of your file. Multi-line
--                  descriptions should align with each other
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:
-- History:
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.registers_pack.all;

entity reg_32b is
    port    (
             Clk      : in  std_logic;                      --  Clk Input
             RST      : in  std_logic;                      --  RST Input
             RdCE     : in  std_logic;                      --  RdCE Input
             WrCE     : in  std_logic;                      --  WrCE Input
             DataIn   : in  std_logic_vector(0 to 31);      --  DataIn Input
             DataOut  : out std_logic_vector(0 to 31);      --  DataOut Output
             RegData  : out std_logic_vector(0 to 31);      --  RegData Output
             TPReq    : out std_logic                       --  TPReq Output
            );
end reg_32b;

------------------------------------------------------------------------------
-- Architecture
------------------------------------------------------------------------------

architecture imp of reg_32b is

------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

signal reg_data : std_logic_vector(0 to 31);
signal wrCE_d   : std_logic;

begin

------------------------------------------------------------------------------
-- Concurrent Signal Assignments
------------------------------------------------------------------------------

RegData   <= reg_data;

------------------------------------------------------------------------------
-- BUS_READ_PROCESS
------------------------------------------------------------------------------

BUS_READ_PROCESS : process (RdCE, reg_data)
begin
    for i in 0 to 31
    loop
        DataOut(i) <= RdCE and reg_data(i);
    end loop;
end process;

------------------------------------------------------------------------------
-- BUS_WRITE_PROCESS
------------------------------------------------------------------------------

BUS_WRITE_PROCESS : process (Clk)
begin
    if (Clk'event and Clk = '1') then
      if (Rst = '1') then
        reg_data <= (others => '0');
        TPReq    <= '0';
        wrCE_d   <= '0';
      elsif (WrCE = '1') then
        reg_data <= DataIn;
        TPReq    <= wrCE_d;
        wrCE_d   <= WrCE;
      else
        TPReq    <= wrCE_d;
        wrCE_d   <= WrCE;
      end if;
    end if;
end process;

end imp;


------------------------------------------------------------------------------
-- $Id: reg_16bl.vhd,v 1.1.2.2 2010/12/15 22:53:05 mwelter Exp $
------------------------------------------------------------------------------
-- reg_16bl - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        reg_16bl.vhd
-- Version:         v2.00a
-- Description:     Include a meaningful description of your file. Multi-line
--                  descriptions should align with each other
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:
-- History:
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.registers_pack.all;

entity reg_16bl is
    port    (
             Clk      : in  std_logic;                      --  Clk Input
             RST      : in  std_logic;                      --  RST Input
             RdCE     : in  std_logic;                      --  RdCE Input
             WrCE     : in  std_logic;                      --  WrCE Input
             DataIn   : in  std_logic_vector(16 to 31);     --  DataIn Input
             DataOut  : out std_logic_vector(16 to 31);     --  DataOut Output
             RegData  : out std_logic_vector(16 to 31);     --  RegData Output
             TPReq    : out std_logic                       --  TPReq Output
            );
end reg_16bl;

------------------------------------------------------------------------------
-- Architecture
------------------------------------------------------------------------------

architecture imp of reg_16bl is

------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------

signal reg_data : std_logic_vector(16 to 31);
signal wrCE_d   : std_logic;

begin

------------------------------------------------------------------------------
-- Concurrent Signal Assignments
------------------------------------------------------------------------------

RegData   <= reg_data;

------------------------------------------------------------------------------
-- BUS_READ_PROCESS
------------------------------------------------------------------------------

BUS_READ_PROCESS : process (RdCE, reg_data)
begin
    for i in 16 to 31
    loop
        DataOut(i) <= RdCE and reg_data(i);
    end loop;
end process;

------------------------------------------------------------------------------
-- BUS_WRITE_PROCESS
------------------------------------------------------------------------------

BUS_WRITE_PROCESS : process (Clk)
begin
    if (Clk'event and Clk = '1') then
      if (Rst = '1') then
        reg_data <= (others => '0');
        TPReq    <= '0';
        wrCE_d   <= '0';
      elsif (WrCE = '1') then
        reg_data <= DataIn;
        TPReq    <= wrCE_d;
        wrCE_d   <= WrCE;
      else
        TPReq    <= wrCE_d;
        wrCE_d   <= WrCE;
      end if;
    end if;
end process;

end imp;


-------------------------------------------------------------------------------
-- reset_combiner - entity/architecture pair
-------------------------------------------------------------------------------
--
-- ***************************************************************************
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of
-- Xilinx, Inc. ("Xilinx"), that is distributed under a license
-- from Xilinx, and may be used, copied and/or disclosed only
-- pursuant to the terms of a valid license agreement with Xilinx.
--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will
-- meet the requirements of Licensee, or that the operation of the
-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2009 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
-- ***************************************************************************
--
-------------------------------------------------------------------------------
-- Filename:        reset_combiner.vhd
-- Version:         v1.00a
-- Description:     combine all resets and capture on proper clock domains
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_uartlite.
--
--              axi_ethernet.vhd
--                reset_combiner.vhd
-------------------------------------------------------------------------------
-- Author:          MSH & MW
--
--  MSH & MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.clock_cross_pack.all;

-------------------------------------------------------------------------------
-- Definition of Generics :
-------------------------------------------------------------------------------
--
--
-------------------------------------------------------------------------------
-- Definition of Ports :
-------------------------------------------------------------------------------
--Inputs
-- BUS2IP_CLK            -- AXI Clock
-- S_AXI_ARESETN         -- AXI Reset
-- Axi_Str_TxD_AClk     --
-- Axi_Str_TxD_AReset   --
-- Axi_Str_TxC_AClk     --
-- Axi_Str_TxC_AReset   --
-- Axi_Str_RxD_AClk     --
-- Axi_Str_rxD_AReset   --
-- Axi_Str_RxS_AClk     --
-- Axi_Str_RxS_AReset   --
--Outputs
-- RESET2AXI
-- saxiResetToAxiStrTxD     --
-- saxiResetToAxiStrTxC     --
-- saxiResetToAxiStrRxD     --
-- saxiResetToAxiStrRxS     --
-------------------------------------------------------------------------------

entity reset_combiner is
    generic (
    C_PHY_RST_COUNT      : integer              := 1321;
    C_FAMILY             : string               := "virtex7";
    C_SIMULATION         : integer range 0 to 1 := 0
);
port (
    S_AXI_ACLK           : in  std_logic;   --  AXI4-Lite Clock
    S_AXI_ARESETN        : in  std_logic;   --  AXI4-Lite Reset
    GTX_CLK_125MHZ       : in  std_logic;   --  GTX CLK
    RX_CLIENT_CLK        : in  std_logic;   --  Receive Client Clock
    RX_CLIENT_CLK_EN     : in  std_logic;   --  Receive Client Clock Enable
    TX_CLIENT_CLK        : in  std_logic;   --  Transmit Client Clock
    TX_CLIENT_CLK_EN     : in  std_logic;   --  Transmit Client Clock Enable
    AXI_STR_TXD_ACLK     : in  std_logic;   --  AXI-Stream Transmit Clock
    AXI_STR_TXD_ARESETN  : in  std_logic;   --  AXI-Stream Transmit Reset
    AXI_STR_TXC_ACLK     : in  std_logic;   --  AXI-Stream Transmit Clock
    AXI_STR_TXC_ARESETN  : in  std_logic;   --  AXI-Stream Transmit Reset
    AXI_STR_RXD_ACLK     : in  std_logic;   --  AXI-Stream Receive Clock
    AXI_STR_RXD_ARESETN  : in  std_logic;   --  AXI-Stream Receive Reset
    AXI_STR_RXS_ACLK     : in  std_logic;   --  AXI-Stream Receive Clock
    AXI_STR_RXS_ARESETN  : in  std_logic;   --  AXI-Stream Receive Reset
    PHY_RESET_N          : out std_logic;   --  PHY Reset
    PHY_RESET_CMPLTE     : out std_logic;   --  PHY Reset Complete
    RESET2AXI            : out std_logic;   --  Reset going to AXI
    RESET2RX_CLIENT      : out std_logic;   --  Reset going to Receive Client Interface
    RESET2TX_CLIENT      : out std_logic;   --  Reset going to Transmit Client Interface
    RESET2AXI_STR_TXD    : out std_logic;   --  Reset going to AXI-Stream Transmit Data Interface
    RESET2AXI_STR_TXC    : out std_logic;   --  Reset going to AXI-Stream Transmit Control Interface
    RESET2AXI_STR_RXD    : out std_logic;   --  Reset going to AXI-Stream Receive Data Interface
    RESET2AXI_STR_RXS    : out std_logic;   --  Reset going to AXI-Stream Receive Status Interface
    RESET2GTX_CLK        : out std_logic    --  Reset going to GTX Clock signals
);
end reset_combiner;

architecture imp of reset_combiner is

    constant C_10MS : unsigned(11 downto 0) := "100000000000"; -- 0x0800
    constant C_15MS : unsigned(11 downto 0) := "110000000000"; -- 0x0C00
    constant C_10US : unsigned(11 downto 0) := "000000000000"; -- 0x01
    constant C_15US : unsigned(11 downto 0) := "000000000001"; -- 0x02

    signal axiStrTxdResetSaxiDomain      : std_logic;
    signal axiStrTxcResetSaxiDomain      : std_logic;
    signal axiStrRxdResetSaxiDomain      : std_logic;
    signal axiStrRxSResetSaxiDomain      : std_logic;

    signal saxiResetAxiStrTxdDomain      : std_logic;
    signal axiStrTxcResetAxiStrTxdDomain : std_logic;
    signal axiStrRxdResetAxiStrTxdDomain : std_logic;
    signal axiStrRxsResetAxiStrTxdDomain : std_logic;

    signal saxiResetAxiStrTxcDomain      : std_logic;
    signal axiStrTxdResetAxiStrTxcDomain : std_logic;
    signal axiStrRxdResetAxiStrTxcDomain : std_logic;
    signal axiStrRxsResetAxiStrTxcDomain : std_logic;

    signal saxiResetAxiStrRxdDomain      : std_logic;
    signal axiStrTxdResetAxiStrRxdDomain : std_logic;
    signal axiStrTxcResetAxiStrRxdDomain : std_logic;
    signal axiStrRxsResetAxiStrRxdDomain : std_logic;

    signal saxiResetAxiStrRxsDomain      : std_logic;
    signal axiStrTxdResetAxiStrRxsDomain : std_logic;
    signal axiStrTxcResetAxiStrRxsDomain : std_logic;
    signal axiStrRxdResetAxiStrRxsDomain : std_logic;

    signal saxiResetGtxDomain            : std_logic;
    signal reset2gtx                     : std_logic;

    signal phy_reset_count               : unsigned(11 downto 0);
    signal reset_delay                   : unsigned(11 downto 0);
    signal reset_done_delay              : unsigned(11 downto 0);

    signal reset2axi_i                   : std_logic;
    signal s_axi_areset                  : std_logic;
    signal axi_str_txd_areset            : std_logic;
    signal axi_str_txc_areset            : std_logic;
    signal axi_str_rxd_areset            : std_logic;
    signal axi_str_rxs_areset            : std_logic;

    signal srl32_1_output                : std_logic;
    signal srl32_2_output                : std_logic;
    signal srl32_2_output_d1             : std_logic;
    signal phyResetCntEnable             : std_logic;

    signal srl32_1_reg                : std_logic_vector (30 downto 0); -- depth is 31
    signal srl32_2_reg                : std_logic_vector (18 downto 0); -- depth is 19

begin

    s_axi_areset       <= not(S_AXI_ARESETN);
    axi_str_txd_areset <= not(AXI_STR_TXD_ARESETN);
    axi_str_txc_areset <= not(AXI_STR_TXC_ARESETN);
    axi_str_rxd_areset <= not(AXI_STR_RXD_ARESETN);
    axi_str_rxs_areset <= not(AXI_STR_RXS_ARESETN);

    NORMAL_DELAY: if(C_SIMULATION = 0) generate
    BEGIN
        reset_delay      <= C_10MS;
        reset_done_delay <= C_15MS;
    end generate NORMAL_DELAY;

    SIMULATION_DELAY: if(C_SIMULATION = 1) generate
    BEGIN
        reset_delay      <= C_10US;
        reset_done_delay <= C_15US;
    end generate SIMULATION_DELAY;


    GEN_UScale: if ( not((C_FAMILY = "kintex7") or (C_FAMILY = "virtex7") or (C_FAMILY = "artix7") or (C_FAMILY = "zynq")))  generate
        PHY_RESET_PULSE : process (S_AXI_ACLK)
        begin
            if (S_AXI_ACLK'event and S_AXI_ACLK = '1') then
                if (s_axi_areset = '1') then
                    phy_reset_count  <= (others => '0');

                    srl32_1_reg <= std_logic_vector(to_unsigned(C_PHY_RST_COUNT,31));
                    if (C_SIMULATION = 1) then
                        srl32_2_reg <= std_logic_vector(to_unsigned(1,19));
                    else 
                        srl32_2_reg <= std_logic_vector(to_unsigned(1000,19));
                    end if ;

                    PHY_RESET_N      <= '0';
                    PHY_RESET_CMPLTE <= '0';
                else
                    if ( phy_reset_count >= 3 ) then
                        srl32_1_reg <= srl32_1_reg;
                    elsif ( unsigned(srl32_1_reg) = 0) then
                        srl32_1_reg <= std_logic_vector(to_unsigned(C_PHY_RST_COUNT,31));
                    else 
                        srl32_1_reg <= std_logic_vector(unsigned(srl32_1_reg) - 1);
                    end if ;

                    if ( ( unsigned(srl32_1_reg) = 0) and (phy_reset_count < 3) ) then
                        if ( unsigned(srl32_2_reg) = 0) then
                            if (C_SIMULATION = 1) then
                                srl32_2_reg <= std_logic_vector(to_unsigned(1,19));
                            else 
                                srl32_2_reg <= std_logic_vector(to_unsigned(1000,19));
                            end if ;
                        else 
                            srl32_2_reg <= std_logic_vector(unsigned(srl32_2_reg) - 1);
                        end if ;
                    else 
                        srl32_2_reg <= srl32_2_reg;
                    end if ;

                    if ( (unsigned(srl32_1_reg) = 0) and (unsigned(srl32_2_reg) = 0) and (phy_reset_count < 3) ) then
                        phy_reset_count <= phy_reset_count + "1";
                    else 
                        phy_reset_count <= phy_reset_count;
                    end if;

                    if ( phy_reset_count < 2 ) then
                        PHY_RESET_N <= '0';
                    else 
                        PHY_RESET_N <= '1';
                    end if;

                    if ( phy_reset_count < 3 ) then
                        PHY_RESET_CMPLTE <= '0';
                    else 
                        PHY_RESET_CMPLTE <= '1';
                    end if;
                end if;
            end if;
        end process;
    end generate GEN_UScale;                                                                           

    GEN_NonUScale: if ((C_FAMILY = "kintex7") or (C_FAMILY = "virtex7") or (C_FAMILY = "artix7") or (C_FAMILY = "zynq"))  generate
        GTX_RESET_PULSE : process (GTX_CLK_125MHZ)
        begin
            if (GTX_CLK_125MHZ'event and GTX_CLK_125MHZ = '1') then
                if (saxiResetGtxDomain = '1') then
                    srl32_2_output_d1        <= '0';
                    phyResetCntEnable        <= '0';
                else
                    srl32_2_output_d1        <= srl32_2_output;
                    phyResetCntEnable        <= srl32_2_output and not(srl32_2_output_d1);
                end if;
            end if;
        end process;

        SRLC32E_1 : process(GTX_CLK_125MHZ)
        begin
            if (GTX_CLK_125MHZ'event and GTX_CLK_125MHZ = '1') then
                if (saxiResetGtxDomain = '1') then      
                    srl32_1_reg <= "0000000000000000000000000000001";
                else
                    srl32_1_reg <= srl32_1_reg(29 downto 0) & srl32_1_reg(30);
                end if;
            end if;
        end process;

        SRLC32E_2 : process(GTX_CLK_125MHZ)
        begin
            if (GTX_CLK_125MHZ'event and GTX_CLK_125MHZ = '1') then
                if (saxiResetGtxDomain = '1') then                 
                    srl32_2_reg <= "0000000000000000001";
                elsif(srl32_1_reg(30)='1') then
                    srl32_2_reg <= srl32_2_reg(17 downto 0) & srl32_2_reg(18);
                end if;
            end if;
        end process;

        srl32_2_output <= srl32_2_reg(18);
  -----------------------------------------------------------------------------
  -- we must hold the PHY reset active for at least 5mS which we will do by
  -- using the known 125 MHz GTX clock
  -----------------------------------------------------------------------------

        COUNT_GTX : process (GTX_CLK_125MHZ)
        begin
            if (GTX_CLK_125MHZ'event and GTX_CLK_125MHZ = '1') then
                if (reset2gtx = '1') then
                    PHY_RESET_N      <= '0';
                    PHY_RESET_CMPLTE <= '0';
                    phy_reset_count  <= (others => '0');
                elsif (phyResetCntEnable = '1') then -- once every 5 uS
                    if (phy_reset_count <= reset_delay) then -- 10mS (10 uS in simulation mode)
                        PHY_RESET_N      <= '0';
                        PHY_RESET_CMPLTE <= '0';
                        phy_reset_count  <= phy_reset_count + 1;
                    elsif (phy_reset_count <= reset_done_delay) then -- 15mS (15 uS in simulation mode)
                        PHY_RESET_N      <= '1';
                        PHY_RESET_CMPLTE <= '0';
                        phy_reset_count  <= phy_reset_count + 1;
                    else
                        PHY_RESET_N  <= '1';
                        PHY_RESET_CMPLTE <= '1';
                    end if;
                end if;
            end if;
        end process;

    end generate GEN_NonUScale;                                                                           


    reset2axi_i      <= s_axi_areset                  or axiStrTxdResetSaxiDomain
                        or axiStrTxcResetSaxiDomain      or axiStrRxdResetSaxiDomain
                        or axiStrRxSResetSaxiDomain;

    RESET2AXI        <= reset2axi_i;

    RESET2AXI_STR_TXD <= saxiResetAxiStrTxdDomain      or axi_str_txd_areset
                         or axiStrTxcResetAxiStrTxdDomain or axiStrRxdResetAxiStrTxdDomain
                         or axiStrRxsResetAxiStrTxdDomain;

    RESET2AXI_STR_TXC <= saxiResetAxiStrTxcDomain      or axiStrTxdResetAxiStrTxcDomain
                         or axi_str_txc_areset            or axiStrRxdResetAxiStrTxcDomain
                         or axiStrRxsResetAxiStrTxcDomain;

    RESET2AXI_STR_RXD <= saxiResetAxiStrRxdDomain      or axiStrTxdResetAxiStrRxdDomain
                         or axiStrTxcResetAxiStrRxdDomain or axi_str_rxd_areset
                         or axiStrRxsResetAxiStrRxdDomain;

    RESET2AXI_STR_RXS <= saxiResetAxiStrRxsDomain      or axiStrTxdResetAxiStrRxsDomain
                         or axiStrTxcResetAxiStrRxsDomain or axiStrRxdResetAxiStrRxsDomain
                         or axi_str_rxs_areset;

    reset2gtx         <= saxiResetGtxDomain;
    RESET2GTX_CLK     <= saxiResetGtxDomain;

    AXI_RESET_TO_RXCLIENT : actv_hi_reset_clk_cross
    port map    (
        ClkA               => S_AXI_ACLK,
        ClkAEN             => '1',
        ClkARst            => reset2axi_i,
        ClkAOutOfClkBRst   => open,
        ClkACombinedRstOut => open,
        ClkB               => RX_CLIENT_CLK,
        ClkBEN             => RX_CLIENT_CLK_EN,
        ClkBRst            => '0',
        ClkBOutOfClkARst   => RESET2RX_CLIENT,
        ClkBCombinedRstOut => open
    );

    AXI_RESET_TO_TXCLIENT : actv_hi_reset_clk_cross
    port map    (
        ClkA               => S_AXI_ACLK,
        ClkAEN             => '1',
        ClkARst            => reset2axi_i,
        ClkAOutOfClkBRst   => open,
        ClkACombinedRstOut => open,
        ClkB               => TX_CLIENT_CLK,
        ClkBEN             => TX_CLIENT_CLK_EN,
        ClkBRst            => '0',
        ClkBOutOfClkARst   => RESET2TX_CLIENT,
        ClkBCombinedRstOut => open
    );

    AXI_RESET_TO_GTX : actv_hi_reset_clk_cross
    port map    (
        ClkA               => S_AXI_ACLK,
        ClkAEN             => '1',
        ClkARst            => s_axi_areset,
        ClkAOutOfClkBRst   => open,
        ClkACombinedRstOut => open,
        ClkB               => GTX_CLK_125MHZ,
        ClkBEN             => '1',
        ClkBRst            => '0',
        ClkBOutOfClkARst   => saxiResetGtxDomain,
        ClkBCombinedRstOut => open
    );

  -----------------------------------------------------------------------------
  -- AXI Reset in
  -----------------------------------------------------------------------------
    AXI_RESET_TO_TXD_AXSTREAM : actv_hi_reset_clk_cross
    port map    
    (
        ClkA               => S_AXI_ACLK,
        ClkAEN             => '1',
        ClkARst            => s_axi_areset,
        ClkAOutOfClkBRst   => axiStrTxdResetSaxiDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_TxD_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_txd_areset,
        ClkBOutOfClkARst   => saxiResetAxiStrTxdDomain,
        ClkBCombinedRstOut => open
    );

    AXI_RESET_TO_TXC_AXSTREAM : actv_hi_reset_clk_cross
    port map    (
        ClkA               => S_AXI_ACLK,
        ClkAEN             => '1',
        ClkARst            => s_axi_areset,
        ClkAOutOfClkBRst   => axiStrTxcResetSaxiDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_TxC_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_txc_areset,
        ClkBOutOfClkARst   => saxiResetAxiStrTxcDomain,
        ClkBCombinedRstOut => open
    );

    AXI_RESET_TO_RXD_AXSTREAM : actv_hi_reset_clk_cross
    port map    (
        ClkA               => S_AXI_ACLK,
        ClkAEN             => '1',
        ClkARst            => s_axi_areset,
        ClkAOutOfClkBRst   => axiStrRxdResetSaxiDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_RxD_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_rxd_areset,
        ClkBOutOfClkARst   => saxiResetAxiStrRxdDomain,
        ClkBCombinedRstOut => open
    );

    AXI_RESET_TO_RXS_AXSTREAM : actv_hi_reset_clk_cross
    port map    (
        ClkA               => S_AXI_ACLK,
        ClkAEN             => '1',
        ClkARst            => s_axi_areset,
        ClkAOutOfClkBRst   => axiStrRxsResetSaxiDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_RxS_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_rxs_areset,
        ClkBOutOfClkARst   => saxiResetAxiStrRxsDomain,
        ClkBCombinedRstOut => open
    );

  -----------------------------------------------------------------------------
  -- AXI Stream TxD Reset in
  -----------------------------------------------------------------------------
    TXD_AXSTREAM_TO_TXC_AXSTREAM : actv_hi_reset_clk_cross
    port map    (
        ClkA               => Axi_Str_TxD_AClk,
        ClkAEN             => '1',
        ClkARst            => axi_str_txd_areset,
        ClkAOutOfClkBRst   => axiStrTxcResetAxiStrTxdDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_TxC_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_txc_areset,
        ClkBOutOfClkARst   => axiStrTxdResetAxiStrTxcDomain,
        ClkBCombinedRstOut => open
    );
    TXD_AXSTREAM_TO_RXD_AXSTREAM : actv_hi_reset_clk_cross
    port map    (
        ClkA               => Axi_Str_TxD_AClk,
        ClkAEN             => '1',
        ClkARst            => axi_str_txd_areset,
        ClkAOutOfClkBRst   => axiStrRxdResetAxiStrTxdDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_RxD_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_rxd_areset,
        ClkBOutOfClkARst   => axiStrTxdResetAxiStrRxdDomain,
        ClkBCombinedRstOut => open
    );
    TXD_AXSTREAM_TO_RXS_AXSTREAM : actv_hi_reset_clk_cross
    port map    (
        ClkA               => Axi_Str_TxD_AClk,
        ClkAEN             => '1',
        ClkARst            => axi_str_txd_areset,
        ClkAOutOfClkBRst   => axiStrRxsResetAxiStrTxdDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_RxS_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_rxs_areset,
        ClkBOutOfClkARst   => axiStrTxdResetAxiStrRxsDomain,
        ClkBCombinedRstOut => open
    );
  -----------------------------------------------------------------------------
  -- AXI Stream TxC Reset in
  -----------------------------------------------------------------------------
    TXC_AXSTREAM_TO_RXD_AXSTREAM : actv_hi_reset_clk_cross
    port map   (
        ClkA               => Axi_Str_TxC_AClk,
        ClkAEN             => '1',
        ClkARst            => axi_str_txc_areset,
        ClkAOutOfClkBRst   => axiStrRxdResetAxiStrTxcDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_RxD_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_rxd_areset,
        ClkBOutOfClkARst   => axiStrTxcResetAxiStrRxdDomain,
        ClkBCombinedRstOut => open
    );
    TXC_AXSTREAM_TO_RXS_AXSTREAM : actv_hi_reset_clk_cross
    port map  (
        ClkA               => Axi_Str_TxC_AClk,
        ClkAEN             => '1',
        ClkARst            => axi_str_txc_areset,
        ClkAOutOfClkBRst   => axiStrRxsResetAxiStrTxcDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_RxS_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_rxs_areset,
        ClkBOutOfClkARst   => axiStrTxcResetAxiStrRxsDomain,
        ClkBCombinedRstOut => open
    );
  -----------------------------------------------------------------------------
  -- AXI Stream RxD Reset in
  -----------------------------------------------------------------------------
    RXD_AXSTREAM_TO_RXS_AXSTREAM : actv_hi_reset_clk_cross
    port map  (
        ClkA               => Axi_Str_RxD_AClk,
        ClkAEN             => '1',
        ClkARst            => axi_str_rxd_areset,
        ClkAOutOfClkBRst   => axiStrRxsResetAxiStrRxdDomain,
        ClkACombinedRstOut => open,
        ClkB               => Axi_Str_RxS_AClk,
        ClkBEN             => '1',
        ClkBRst            => axi_str_rxs_areset,
        ClkBOutOfClkARst   => axiStrRxdResetAxiStrRxsDomain,
        ClkBCombinedRstOut => open
    );
end imp;


------------------------------------------------------------------------
-- Title      : Package for the tx_if logic
-- Project    : Tri-Mode Ethernet FIFO
------------------------------------------------------------------------
-- File       : tx_if_pack.vhd
-- Author     : Xilinx Inc.
------------------------------------------------------------------------
-- (c) Copyright 2012 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
------------------------------------------------------------------------
-- Description:  This package contains all component declarations for
--               the entiries which make up the Tx I/F logic
------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;



package tx_if_pack is


  component tx_if
  generic (
    C_FAMILY               : string                        := "virtex6";
    C_HALFDUP              : integer range 0 to 1          := 0;
    C_SPEED_2P5            : integer range 0 to 1          := 0;
    C_TXCSUM               : integer range 0 to 2          := 0;
    C_TXMEM                : integer                       := 4096;
    C_ENABLE_1588       : integer   := 0;
    C_TXVLAN_TRAN          : integer range 0 to 1          := 0;
    C_TXVLAN_TAG           : integer range 0 to 1          := 0;
    C_TXVLAN_STRP          : integer range 0 to 1          := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32        := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32        := 32
  );
  port (

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK                 : in  std_logic;                                     --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd                : in  std_logic;                                     --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID               : in  std_logic;                                     --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY               : out std_logic;                                     --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST                : in  std_logic;                                     --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB                : in  std_logic_vector(3 downto 0);                  --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA                : in  std_logic_vector(31 downto 0);                 --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK                 : in  std_logic;                                     --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc                : in  std_logic;                                     --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID               : in  std_logic;                                     --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY               : out std_logic;                                     --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST                : in  std_logic;                                     --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB                : in  std_logic_vector(3 downto 0);                  --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA                : in  std_logic_vector(31 downto 0);                 --  AXI-Stream Transmit Control Data

    -- VLAN Interface
    tx_vlan_bram_addr                : out std_logic_vector(11 downto 0);                 --  Transmit VLAN BRAM Addr
    tx_vlan_bram_din                 : in  std_logic_vector(13 downto 0);                 --  Transmit VLAN BRAM Rd Data
    tx_vlan_bram_en                  : out std_logic;                                     --  Transmit VLAN BRAM Enable

    enable_newFncEn                  : out std_logic; --Only perform VLAN when FLAG = 0xA --  Enable Extended VLAN Functions
    transMode_cross                  : in  std_logic;                                     --  VLAN Translation Mode Control Bit
    tagMode_cross                    : in  std_logic_vector( 1 downto 0);                 --  VLAN TAG Mode Control Bits
    strpMode_cross                   : in  std_logic_vector( 1 downto 0);                 --  VLAN Strip Mode Control Bits

    tpid0_cross                      : in  std_logic_vector(15 downto 0);                 --  VLAN TPID
    tpid1_cross                      : in  std_logic_vector(15 downto 0);                 --  VLAN TPID
    tpid2_cross                      : in  std_logic_vector(15 downto 0);                 --  VLAN TPID
    tpid3_cross                      : in  std_logic_vector(15 downto 0);                 --  VLAN TPID

    newTagData_cross                 : in  std_logic_vector(31 downto 0);                 --  VLAN Tag Data

    tx_init_in_prog                  : out std_logic;                                     --  Tx is Initializing after a reset
    tx_init_in_prog_cross            : in  std_logic;                                     --  Tx is Initializing after a reset



    tx_mac_aclk                      : in  std_logic;                                 --  Tx AXI-Stream clock in
    tx_reset                         : in  std_logic;                                 --  take to reset combiner
    tx_axis_mac_tdata                : out std_logic_vector(7 downto 0);              --  Tx AXI-Stream data
    tx_axis_mac_tvalid               : out std_logic;                                 --  Tx AXI-Stream valid
    tx_axis_mac_tlast                : out std_logic;                                 --  Tx AXI-Stream last
    tx_axis_mac_tuser                : out std_logic;                  -- this is always driven low since an underflow cannot occur
    tx_axis_mac_tready               : in  std_logic;                                 --  Tx AXI-Stream ready in from TEMAC
    tx_collision                     : in  std_logic;                                 --  collision not used
    tx_retransmit                    : in  std_logic;                                 -- retransmit not used

    tx_client_10_100                 : in  std_logic;                                 --  Tx Client CE Toggles Indicator
    tx_cmplt                         : out std_logic                                  -- transmit is complete indicator

  );
  end component;


  component tx_emac_if
  generic (
    C_FAMILY                  : string                      := "virtex6";
    C_HALFDUP                 : integer range 0 to 1        := 0;
    C_TXMEM                   : integer                     := 4096;
    C_TXCSUM                  : integer range 0 to 2        := 0;
    C_ENABLE_1588       : integer   := 0;

    -- Read Port - AXI Stream TxData
    c_TxD_write_width_a       : integer range   0 to 18     := 9;
    c_TxD_read_width_a        : integer range   0 to 18     := 9;
    c_TxD_write_depth_a       : integer range   0 to 32768  := 4096;
    c_TxD_read_depth_a        : integer range   0 to 32768  := 4096;
    c_TxD_addra_width         : integer range   0 to 15     := 10;
    c_TxD_wea_width           : integer range   0 to 2      := 2;

    -- Read Port - AXI Stream TxControl
    c_TxC_write_width_a       : integer range  36 to 36     := 36;
    c_TxC_read_width_a        : integer range  36 to 36     := 36;
    c_TxC_write_depth_a       : integer range   0 to 1024   := 1024;
    c_TxC_read_depth_a        : integer range   0 to 1024   := 1024;
    c_TxC_addra_width         : integer range   0 to 10     := 10;
    c_TxC_wea_width           : integer range   0 to 1      := 1;

    c_TxD_addrb_width         : integer range   0 to 13     := 10;

    C_CLIENT_WIDTH            : integer                     := 8
  );
  port (
    --Transmit Memory Read Interface
    tx_client_10_100          : in  std_logic;                                        --  Tx Client CE Toggles Indicator
      -- ** WARNING ** WARNING ** WARNING **
      --  For MII,GMII, RGMI, 1000Base-X and pcs/pma SGMII this is an accurate indicator
      --  However for V6 Hard SGMII it is always tied to '0' for all speeds


    -- Read Port - AXI Stream TxData
    reset2tx_client           : in  std_logic;                                        --  reset
    Tx_Client_TxD_2_Mem_Din   : out std_logic_vector(c_TxD_write_width_a-1 downto 0); --  Tx AXI-Stream Data to Memory Wr Din
    Tx_Client_TxD_2_Mem_Addr  : out std_logic_vector(c_TxD_addra_width-1   downto 0); --  Tx AXI-Stream Data to Memory Wr Addr
    Tx_Client_TxD_2_Mem_En    : out std_logic;                                        --  Tx AXI-Stream Data to Memory Enable
    Tx_Client_TxD_2_Mem_We    : out std_logic_vector(c_TxD_wea_width-1     downto 0); --  Tx AXI-Stream Data to Memory Wr En
    Tx_Client_TxD_2_Mem_Dout  : in  std_logic_vector(c_TxD_read_width_a-1  downto 0); --  Tx AXI-Stream Data to Memory Not Used

    -- Read Port - AXI Stream TxControl
    reset2axi_str_txd         : in  std_logic;                                        --  reset
    Tx_Client_TxC_2_Mem_Din   : out std_logic_vector(c_TxC_write_width_a-1 downto 0); --  Tx AXI-Stream Control to Memory Wr Din
    Tx_Client_TxC_2_Mem_Addr  : out std_logic_vector(c_TxC_addra_width-1   downto 0); --  Tx AXI-Stream Control to Memory Wr Addr
    Tx_Client_TxC_2_Mem_En    : out std_logic;                                        --  Tx AXI-Stream Control to Memory Enable
    Tx_Client_TxC_2_Mem_We    : out std_logic_vector(c_TxC_wea_width-1     downto 0); --  Tx AXI-Stream Control to Memory Wr En
    Tx_Client_TxC_2_Mem_Dout  : in  std_logic_vector(c_TxC_read_width_a-1  downto 0); --  Tx AXI-Stream Control to Memory Full Flag

    --  Tx AXI-S Interface
    tx_axi_clk                : in  std_logic;                                        --  Tx AXI-Stream clock in
    tx_reset_out              : in  std_logic;                                        --  take to reset combiner
    tx_axis_mac_tdata         : out std_logic_vector(C_CLIENT_WIDTH - 1 downto 0);    --  Tx AXI-Stream data
    tx_axis_mac_tvalid        : out std_logic;                                        --  Tx AXI-Stream valid
    tx_axis_mac_tlast         : out std_logic;                                        --  Tx AXI-Stream last
    tx_axis_mac_tuser         : out std_logic;                         -- this is always driven low since an underflow cannot occur
    tx_axis_mac_tready        : in  std_logic;                                        --  Tx AXI-Stream ready in from TEMAC
    tx_collision              : in  std_logic;                                        --  collision not used
    tx_retransmit             : in  std_logic;                                        -- retransmit not used


    tx_cmplt                  : out std_logic;                                        -- transmit is complete indicator

    tx_init_in_prog_cross     : in  std_logic                                         --  Tx is Initializing after a reset
  );
  end component;
  
  component tx_emac_if_2g5
  generic (
    C_FAMILY                  : string                      := "virtex6";
    C_HALFDUP                 : integer range 0 to 1        := 0;
    C_TXMEM                   : integer                     := 4096;
    C_TXCSUM                  : integer range 0 to 2        := 0;
    C_ENABLE_1588       : integer   := 0;

    -- Read Port - AXI Stream TxData
    c_TxD_write_width_a       : integer range   0 to 18     := 9;
    c_TxD_read_width_a        : integer range   0 to 18     := 9;
    c_TxD_write_depth_a       : integer range   0 to 32768  := 4096;
    c_TxD_read_depth_a        : integer range   0 to 32768  := 4096;
    c_TxD_addra_width         : integer range   0 to 15     := 10;
    c_TxD_wea_width           : integer range   0 to 2      := 2;

    -- Read Port - AXI Stream TxControl
    c_TxC_write_width_a       : integer range  36 to 36     := 36;
    c_TxC_read_width_a        : integer range  36 to 36     := 36;
    c_TxC_write_depth_a       : integer range   0 to 1024   := 1024;
    c_TxC_read_depth_a        : integer range   0 to 1024   := 1024;
    c_TxC_addra_width         : integer range   0 to 10     := 10;
    c_TxC_wea_width           : integer range   0 to 1      := 1;

    c_TxD_addrb_width         : integer range   0 to 13     := 10;

    C_CLIENT_WIDTH            : integer                     := 8
  );
  port (
    --Transmit Memory Read Interface
    tx_client_10_100          : in  std_logic;                                        --  Tx Client CE Toggles Indicator
      -- ** WARNING ** WARNING ** WARNING **
      --  For MII,GMII, RGMI, 1000Base-X and pcs/pma SGMII this is an accurate indicator
      --  However for V6 Hard SGMII it is always tied to '0' for all speeds


    -- Read Port - AXI Stream TxData
    reset2tx_client           : in  std_logic;                                        --  reset
    Tx_Client_TxD_2_Mem_Din   : out std_logic_vector(c_TxD_write_width_a-1 downto 0); --  Tx AXI-Stream Data to Memory Wr Din
    Tx_Client_TxD_2_Mem_Addr  : out std_logic_vector(c_TxD_addra_width-1   downto 0); --  Tx AXI-Stream Data to Memory Wr Addr
    Tx_Client_TxD_2_Mem_En    : out std_logic;                                        --  Tx AXI-Stream Data to Memory Enable
    Tx_Client_TxD_2_Mem_We    : out std_logic_vector(c_TxD_wea_width-1     downto 0); --  Tx AXI-Stream Data to Memory Wr En
    Tx_Client_TxD_2_Mem_Dout  : in  std_logic_vector(c_TxD_read_width_a-1  downto 0); --  Tx AXI-Stream Data to Memory Not Used

    -- Read Port - AXI Stream TxControl
    reset2axi_str_txd         : in  std_logic;                                        --  reset
    Tx_Client_TxC_2_Mem_Din   : out std_logic_vector(c_TxC_write_width_a-1 downto 0); --  Tx AXI-Stream Control to Memory Wr Din
    Tx_Client_TxC_2_Mem_Addr  : out std_logic_vector(c_TxC_addra_width-1   downto 0); --  Tx AXI-Stream Control to Memory Wr Addr
    Tx_Client_TxC_2_Mem_En    : out std_logic;                                        --  Tx AXI-Stream Control to Memory Enable
    Tx_Client_TxC_2_Mem_We    : out std_logic_vector(c_TxC_wea_width-1     downto 0); --  Tx AXI-Stream Control to Memory Wr En
    Tx_Client_TxC_2_Mem_Dout  : in  std_logic_vector(c_TxC_read_width_a-1  downto 0); --  Tx AXI-Stream Control to Memory Full Flag

    --  Tx AXI-S Interface
    tx_axi_clk                : in  std_logic;                                        --  Tx AXI-Stream clock in
    tx_reset_out              : in  std_logic;                                        --  take to reset combiner
    tx_axis_mac_tdata         : out std_logic_vector(C_CLIENT_WIDTH - 1 downto 0);    --  Tx AXI-Stream data
    tx_axis_mac_tvalid        : out std_logic;                                        --  Tx AXI-Stream valid
    tx_axis_mac_tlast         : out std_logic;                                        --  Tx AXI-Stream last
    tx_axis_mac_tuser         : out std_logic;                         -- this is always driven low since an underflow cannot occur
    tx_axis_mac_tready        : in  std_logic;                                        --  Tx AXI-Stream ready in from TEMAC
    tx_collision              : in  std_logic;                                        --  collision not used
    tx_retransmit             : in  std_logic;                                        -- retransmit not used


    tx_cmplt                  : out std_logic;                                        -- transmit is complete indicator

    tx_init_in_prog_cross     : in  std_logic                                         --  Tx is Initializing after a reset
  );
  end component;


  component tx_csum_partial_if
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data


    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0)   --  Tx AXI-Stream Control to Memory Full Flag

  );
  end component;


  component tx_csum_partial_calc_if
  generic (
    C_FAMILY                  : string                      := "virtex6";
    C_TXCSUM                  : integer range 0 to 2        := 0;
    C_S_AXI_DATA_WIDTH        : integer range 32 to 32      := 32;
    c_TxD_addrb_width         : integer range  0 to 13      := 10
  );
  port (
    AXI_STR_TXC_ACLK           : in  std_logic;                                       --  AXI-Stream Transmit Control Clock
    reset2axi_str_txc          : in  std_logic;                                       --  Reset
    axi_str_txc_tready_int_dly : in  std_logic;                                       --  AXI-Stream Transmit Control Ready
    axi_str_txc_tvalid_dly0    : in  std_logic;                                       --  AXI-Stream Transmit Control Valid
    axi_str_txc_tlast_dly0     : in  std_logic;                                       --  AXI-Stream Transmit Control Last

    load_csum_int              : in  std_logic;                                       --  Load CSUM Initial Value
    axi_flag                   : in  std_logic_vector( 3 downto 0);                   --  AXI Flag From AXI-Stream Tx Control
    csum_cntrl                 : in  std_logic_vector( 1 downto 0);                   --  CSUM Control Bits = "01" for partial CSUM
    csum_begin                 : in  std_logic_vector(c_TxD_addrb_width -1 downto 0); --  CSUM Start Location
    csum_begin_bytes           : in  std_logic_vector( 1 downto 0);                   --  CSUM Enables for which Byte to start calc
    csum_insert                : in  std_logic_vector(c_TxD_addrb_width -1 downto 0); --  CSUM Insertion Location
    csum_insert_bytes          : in  std_logic_vector( 1 downto 0);                   --  CSUM Enables for which Byte to insert at
    csum_init                  : in  std_logic_vector(15 downto 0);                   --  CSUM INitial Value to start at

    AXI_STR_TXD_ACLK           : in  std_logic;                                       --  AXI-Stream Transmit Data Clock
    reset2axi_str_txd          : in  std_logic;                                       --  Reset
    csum_addr                  : in  std_logic_vector(c_TxD_addrb_width -1 downto 0); --  Current address to Tx Data Memory
    inc_txd_wr_addr            : in  std_logic;                                       --  Incraments the Wr address
    inc_txd_addr_one           : in  std_logic;                                       --  Incraments the Wr address at the end
    non_xilinx_ip_pulse        : in  std_logic;                                       --  Not Supported
    axi_str_txd_tdata_dly1     : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0); --  AXI-Stream Transmit Memory Data

    do_csum                    : out std_logic;                                       --  Enable to do CSUM
    csum_result                : out std_logic_vector(15 downto 0);                   --  Final CSUM result valid with csum_en
    csum_en                    : out std_logic;                                       --  Final CSUM resullt is valid
    csum_we                    : out std_logic_vector(3 downto 0);                    --  Memory Write Enables for 16-bit access
    csum_cmplt                 : out std_logic                                        --  Current CSUM calculation is complete
  );

  end component;


  component tx_csum_if
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0)   --  Tx AXI-Stream Control to Memory Full Flag

  );

  end component;


  component tx_csum_full_if
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data


    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0)   --  Tx AXI-Stream Control to Memory Full Flag

  );
  end component;


  component tx_csum_full_fsm
  generic (
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32     := 32;
    c_TxD_addrb_width      : integer range  0 to 13     := 10
  );
  port (

    AXI_STR_TXD_ACLK  : in  std_logic;                                        --  Clock
    reset2axi_str_txd : in  std_logic;                                        --  Reset

    txd_strbs         : in  std_logic_vector(3 downto 0);                     --  AXI-Stream Tx Data Strobes
    do_csum           : in  std_logic;                                        --  axi_flag must = 0xA for this to be enabled
    abort_csum        : out std_logic;                                        --  All conditions were not met to complete csum
    txd_tlast         : in  std_logic;                                        --  AXI-Stream Tx Data Last
    csum_calc_en      : in  std_logic;                                        --  axi_str_txd_tvalid_dly0 and
                                                                              --  axi_str_txd_tready_int_dly;
    clr_csums         : out std_logic;                                        --  Clear CSUM flags and calculations
    tcp_ptcl          : out std_logic;                                        --  TCP Protocol Indicator
    udp_ptcl          : out std_logic;                                        --  UDP Protocol Indicator
    en_ipv4_hdr_b32   : out std_logic_vector( 1 downto 0);                    --  bytes 3 and 2 of din
    en_ipv4_hdr_b10   : out std_logic_vector( 1 downto 0);                    --  bytes 1 and 0 of din
    last_ipv4_hdr_cnt : out std_logic;                                        --  last data for IPv4 Header Calculation
    fsm_csum_en_b32   : out std_logic_vector( 1 downto 0);                    --  bytes 3 and 2 of din
    fsm_csum_en_b10   : out std_logic_vector( 1 downto 0);                    --  bytes 1 and 0 of din
    add_psdo_wd       : out std_logic;                                        --  last data for TCP/UDP Calculation
    ptcl_csum_cmplt   : in  std_logic;                                        --  indicates the TCP/UDP csum calculation is complete
    zeroes_en         : out std_logic_vector( 1 downto 0);                    --  stalls the CSUM calculations for one clock so
                                                                              --  Zeroes do not need muxed in
    din               : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1  downto 0); --  AXI Stream Tx Data
    csum_din          : out std_logic_vector(C_S_AXI_DATA_WIDTH-1  downto 0); --  Mux out of pseudo data or axi_str_txd_tdata_dly0
    do_ipv4hdr        : out std_logic;                                        --  only do the ipv4 header csum
    not_tcp_udp       : out std_logic;                                        --  only do the ipv4 header csum - no TCP/UDP protocol
    do_full_csum      : out std_logic;                                        --  do the ipv4 headr and TCP/UDP csum
    hdr_csum_cmplt    : in  std_logic;                                        --  Header CSUM Calculation is complete
    wr_hdr_csum       : out std_logic;                                        --  Enable to Write the Header CSUM to Memory
    wr_ptcl_csum      : out std_logic;                                        --  Enable to Write the EthII/Snap Ipv4 TCP/UDP CSUM

    csum_strt_addr    : in  std_logic_vector(c_TxD_addrb_width-1   downto 0); --  Start Address to start the CSUM ccalculation
    csum_ipv4_hdr_addr: out std_logic_vector(c_TxD_addrb_width-1   downto 0); --  IPv4 Header Start Address
    csum_ipv4_hdr_we  : out std_logic_vector( 3 downto 0);                    --  IPv4 Header Write Enable to Memory
    csum_ptcl_addr    : out std_logic_vector(c_TxD_addrb_width-1   downto 0); --  Address to Write the EthII/Snap Ipv4 TCP/UDP CSUM
    csum_ptcl_we      : out std_logic_vector( 3 downto 0)                     --  Enables to Write the EthII/Snap Ipv4 TCP/UDP CSUM
  );
  end component;


  component tx_csum_full_calc_if
  generic (
    -- 0 = calculate the TCP/UDP CSUM
    -- 1 = calculate the IPv4 Header CSUM
    C_IPV4_HEADER_CSUM  : integer range 0 to 1 := 0
  );
  port (
    clk               : in  std_logic;                      --  clk
    reset             : in  std_logic;                      --  reset
    clr_csums         : in  std_logic;                      --  clear the csum
    txd_tlast         : in  std_logic;                      --  axi_str_txd_tlast_dly0,
    csum_calc_en      : in  std_logic;                      --  axi_str_txd_tvalid_dly0 and axi_str_txd_tready_int_dly;

    tcp_ptcl          : in  std_logic;                      --  tcp protocol flag
    udp_ptcl          : in  std_logic;                      --  udp protocol flag
    do_ipv4hdr        : in  std_logic;                      --  only do the ipv4 header csum
    not_tcp_udp       : in  std_logic;                      --  only do the ipv4 header csum after received tlast in ptcol header
    do_full_csum      : in  std_logic;                      --  do IPv4 Ethernet II or SNAP CSUM

    do_csum           : in  std_logic;                      --  Full CSUM FLAG is set
    csum_en_b32       : in  std_logic_vector(1 downto 0);   --  enables for either IPv4 header or TCP/UDP CSUM calc bytes 3,2
    csum_en_b10       : in  std_logic_vector(1 downto 0);   --  enables for either IPv4 header or TCP/UDP CSUM calc bytes 1,0
    zeroes_en         : in  std_logic_vector(1 downto 0);   --  zeroes for either IPv4 header or TCP/UDP CSUM calc

    data_last         : in  std_logic;                      --  last data to be included in the csum calculation
    inc_txd_addr_one  : in  std_logic;                       --  increments the Tx Data Memory Address at end of a packet
    inc_txd_addr_one_early : in  std_logic;                 --  Pulses onle clock cycle early when do_csum is enabled with
                                                            --  txd_tlast and csum_calc_en

    csum_din          : in  std_logic_vector(31 downto 0);  --  Data for CSUM calculation
    csum_dout         : out std_logic_vector(15 downto 0);  --  Computed CSUM Result
    csum_we           : out std_logic_vector( 3 downto 0);  --  Tx Data Memory Write Enables to perform 16-bit write
    csum_cmplt        : out std_logic                       --  CSUM Calculation has completed
  );
  end component;

  component  tx_vlan_if 
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_TYPE                 : integer range 0 to 2         := 0;
    C_PHY_TYPE             : integer range 0 to 7         := 1;
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data

    --Transmit EMAC Interface

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0);  --  Tx AXI-Stream Control to Memory Full Flag

    tx_vlan_bram_addr      : out std_logic_vector(11 downto 0);                     --  Transmit VLAN BRAM Addr
    tx_vlan_bram_din       : in  std_logic_vector(13 downto 0);                     --  Transmit VLAN BRAM Rd Data
    tx_vlan_bram_en        : out std_logic;                                         --  Transmit VLAN BRAM Enable

    enable_newFncEn        : out std_logic; --Only perform VLAN when the FLAG = 0xA --  Enable Extended VLAN Functions
    transMode_cross        : in  std_logic;                                         --  VLAN Translation Mode Control Bit
    tagMode_cross          : in  std_logic_vector( 1 downto 0);                     --  VLAN TAG Mode Control Bits
    strpMode_cross         : in  std_logic_vector( 1 downto 0);                     --  VLAN Strip Mode Control Bits

    tpid0_cross            : in  std_logic_vector(15 downto 0);                     --  VLAN TPID
    tpid1_cross            : in  std_logic_vector(15 downto 0);                     --  VLAN TPID
    tpid2_cross            : in  std_logic_vector(15 downto 0);                     --  VLAN TPID
    tpid3_cross            : in  std_logic_vector(15 downto 0);                     --  VLAN TPID

    newTagData_cross       : in  std_logic_vector(31 downto 0)                      --  VLAN Tag Data

  );
  end component;


  component tx_basic_if
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0)   --  Tx AXI-Stream Control to Memory Full Flag

  );
  end component;


  component tx_axistream_if
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                           --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                           --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                           --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                           --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                           --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                        --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);     --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                           --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                           --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                           --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                           --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                           --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                        --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);     --  AXI-Stream Transmit Control Data


    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);    --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);    --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                           --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);    --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);    --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);    --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);    --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                           --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);    --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0);    --  Tx AXI-Stream Control to Memory Full Flag

    -- VLAN Signals
    tx_vlan_bram_addr      : out std_logic_vector(11 downto 0);                       --  Transmit VLAN BRAM Addr
    tx_vlan_bram_din       : in  std_logic_vector(13 downto 0);                       --  Transmit VLAN BRAM Rd Data
    tx_vlan_bram_en        : out std_logic;                                           --  Transmit VLAN BRAM Enable

    enable_newFncEn        : out std_logic; --Only perform VLAN when the FLAG = 0xA   --  Enable Extended VLAN Functions
    transMode_cross        : in  std_logic;                                           --  VLAN Translation Mode Control Bit
    tagMode_cross          : in  std_logic_vector( 1 downto 0);                       --  VLAN TAG Mode Control Bits
    strpMode_cross         : in  std_logic_vector( 1 downto 0);                       --  VLAN Strip Mode Control Bits

    tpid0_cross            : in  std_logic_vector(15 downto 0);                       --  VLAN TPID
    tpid1_cross            : in  std_logic_vector(15 downto 0);                       --  VLAN TPID
    tpid2_cross            : in  std_logic_vector(15 downto 0);                       --  VLAN TPID
    tpid3_cross            : in  std_logic_vector(15 downto 0);                       --  VLAN TPID

    newTagData_cross       : in  std_logic_vector(31 downto 0);                       --  VLAN Tag Data

    tx_init_in_prog        : out std_logic                                            --  Tx is Initializing after a reset

  );
  end component;


  component tx_mem_if
  generic (
    C_FAMILY               : string                      := "virtex6";

    -- Read Port - AXI Stream TxData
    c_TxD_write_width_a      : integer range   0 to 18     := 9;
    c_TxD_read_width_a       : integer range   0 to 18     := 9;
    c_TxD_write_depth_a      : integer range   0 to 32768  := 4096;
    c_TxD_read_depth_a       : integer range   0 to 32768  := 4096;
    c_TxD_addra_width        : integer range   0 to 15     := 10;
    c_TxD_wea_width          : integer range   0 to 2      := 2;
    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b      : integer range  36 to 36     := 36;
    c_TxD_read_width_b       : integer range  36 to 36     := 36;
    c_TxD_write_depth_b      : integer range   0 to 8192   := 1024;
    c_TxD_read_depth_b       : integer range   0 to 8192   := 1024;
    c_TxD_addrb_width        : integer range   0 to 13     := 10;
    c_TxD_web_width          : integer range   0 to 4      := 4;

    -- Read Port - AXI Stream TxControl
    c_TxC_write_width_a      : integer range  36 to 36     := 36;
    c_TxC_read_width_a       : integer range  36 to 36     := 36;
    c_TxC_write_depth_a      : integer range   0 to 1024   := 1024;
    c_TxC_read_depth_a       : integer range   0 to 1024   := 1024;
    c_TxC_addra_width        : integer range   0 to 10     := 10;
    c_TxC_wea_width          : integer range   0 to 1      := 1;
    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b      : integer range   36 to 36    := 36;
    c_TxC_read_width_b       : integer range   36 to 36    := 36;
    c_TxC_write_depth_b      : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b       : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width        : integer range    0 to 10    := 10;
    c_TxC_web_width          : integer range    0 to 1     := 1

  );
  port (
    -- Read Port - AXI Stream TxData
    TX_CLIENT_CLK             : in  std_logic;                                          --  Tx Client Clock
    reset2tx_client           : in  std_logic;                                          --  Reset
    Tx_Client_TxD_2_Mem_Din   : in  std_logic_vector(c_TxD_write_width_a-1 downto 0);   --  Tx Client Data Memory Wr Data
    Tx_Client_TxD_2_Mem_Addr  : in  std_logic_vector(c_TxD_addra_width-1   downto 0);   --  Tx Client Data Memory Address
    Tx_Client_TxD_2_Mem_En    : in  std_logic;                                          --  Tx Client Data Memory Enable
    Tx_Client_TxD_2_Mem_We    : in  std_logic_vector(c_TxD_wea_width-1     downto 0);   --  Tx Client Data Memory Wr Enable
    Tx_Client_TxD_2_Mem_Dout  : out std_logic_vector(c_TxD_read_width_a-1  downto 0);   --  Tx Client Data Memory Rd Data
    -- Write Port - AXI Stream TxData
    AXI_STR_TXD_ACLK          : in  std_logic;                                          --  AXI-Stream Tx Data Clock
    reset2axi_str_txd         : in  std_logic;                                          --  Reset
    Axi_Str_TxD_2_Mem_Din     : in  std_logic_vector(c_TxD_write_width_b-1 downto 0);   --  AXI-Stream Tx Data Memory Wr Data
    Axi_Str_TxD_2_Mem_Addr    : in  std_logic_vector(c_TxD_addrb_width-1   downto 0);   --  AXI-Stream Tx Data Memory Address
    Axi_Str_TxD_2_Mem_En      : in  std_logic;                                          --  AXI-Stream Tx Data Memory Enable
    Axi_Str_TxD_2_Mem_We      : in  std_logic_vector(c_TxD_web_width-1     downto 0);   --  AXI-Stream Tx Data Memory Wr Enable
    Axi_Str_TxD_2_Mem_Dout    : out std_logic_vector(c_TxD_read_width_b-1  downto 0);   --  AXI-Stream Tx Data Memory Rd Data

    -- Read Port - AXI Stream TxControl
    Tx_Client_TxC_2_Mem_Din   : in  std_logic_vector(c_TxC_write_width_a-1 downto 0);   --  Tx Client Control Memory Wr Data
    Tx_Client_TxC_2_Mem_Addr  : in  std_logic_vector(c_TxC_addra_width-1   downto 0);   --  Tx Client Control Memory Address
    Tx_Client_TxC_2_Mem_En    : in  std_logic;                                          --  Tx Client Control Memory Enable
    Tx_Client_TxC_2_Mem_We    : in  std_logic_vector(c_TxC_wea_width-1     downto 0);   --  Tx Client Control Memory Wr Enable
    Tx_Client_TxC_2_Mem_Dout  : out std_logic_vector(c_TxC_read_width_a-1  downto 0);   --  Tx Client Control Memory Rd Data
    -- Write Port - AXI Stream TxControl
    AXI_STR_TXC_ACLK          : in  std_logic;                                          --  AXI-Stream Tx Control Clock
    reset2axi_str_txc         : in  std_logic;                                          --  Reset
    Axi_Str_TxC_2_Mem_Din     : in  std_logic_vector(c_TxC_write_width_b-1 downto 0);   --  AXI-Stream Tx Control Memory Wr Data
    Axi_Str_TxC_2_Mem_Addr    : in  std_logic_vector(c_TxC_addrb_width-1   downto 0);   --  AXI-Stream Tx Control Memory Address
    Axi_Str_TxC_2_Mem_En      : in  std_logic;                                          --  AXI-Stream Tx Control Memory Enable
    Axi_Str_TxC_2_Mem_We      : in  std_logic_vector(c_TxC_web_width-1     downto 0);   --  AXI-Stream Tx Control Memory Wr Enable
    Axi_Str_TxC_2_Mem_Dout    : out std_logic_vector(c_TxC_read_width_b-1  downto 0)    --  AXI-Stream Tx Control Memory Rd Data
  );
  end component;


end tx_if_pack;


-------------------------------------------------------------------------------
-- tx_csum_partial_calc_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_csum_partial_calc_if.vhd
-- Version:         v1.00a
-- Description:     top level of embedded ip Ethernet MAC interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--                    tx_axistream_if.vhd
--                      tx_basic_if.vhd
--                      tx_csum_if.vhd
--                        tx_csum_partial_if.vhd
--          ->              tx_csum_partial_calc_if.vhd
--                        tx_full_csum_if.vhd
--                      tx_vlan_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tx_if_pack.all;


-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity tx_csum_partial_calc_if is
  generic (
    C_FAMILY                  : string                      := "virtex6";
    C_TXCSUM                  : integer range 0 to 2        := 0;
    C_S_AXI_DATA_WIDTH        : integer range 32 to 32      := 32;
    c_TxD_addrb_width         : integer range  0 to 13      := 10
  );
  port (
    AXI_STR_TXC_ACLK           : in  std_logic;                                       --  AXI-Stream Transmit Control Clock
    reset2axi_str_txc          : in  std_logic;                                       --  Reset
    axi_str_txc_tready_int_dly : in  std_logic;                                       --  AXI-Stream Transmit Control Ready
    axi_str_txc_tvalid_dly0    : in  std_logic;                                       --  AXI-Stream Transmit Control Valid
    axi_str_txc_tlast_dly0     : in  std_logic;                                       --  AXI-Stream Transmit Control Last

    load_csum_int              : in  std_logic;                                       --  Load CSUM Initial Value
    axi_flag                   : in  std_logic_vector( 3 downto 0);                   --  AXI Flag From AXI-Stream Tx Control
    csum_cntrl                 : in  std_logic_vector( 1 downto 0);                   --  CSUM Control Bits = "01" for partial CSUM
    csum_begin                 : in  std_logic_vector(c_TxD_addrb_width -1 downto 0); --  CSUM Start Location
    csum_begin_bytes           : in  std_logic_vector( 1 downto 0);                   --  CSUM Enables for which Byte to start calc
    csum_insert                : in  std_logic_vector(c_TxD_addrb_width -1 downto 0); --  CSUM Insertion Location
    csum_insert_bytes          : in  std_logic_vector( 1 downto 0);                   --  CSUM Enables for which Byte to insert at
    csum_init                  : in  std_logic_vector(15 downto 0);                   --  CSUM INitial Value to start at

    AXI_STR_TXD_ACLK           : in  std_logic;                                       --  AXI-Stream Transmit Data Clock
    reset2axi_str_txd          : in  std_logic;                                       --  Reset
    csum_addr                  : in  std_logic_vector(c_TxD_addrb_width -1 downto 0); --  Current address to Tx Data Memory
    inc_txd_wr_addr            : in  std_logic;                                       --  Incraments the Wr address
    inc_txd_addr_one           : in  std_logic;                                       --  Incraments the Wr address at the end
    non_xilinx_ip_pulse        : in  std_logic;                                       --  Not Supported
    axi_str_txd_tdata_dly1     : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0); --  AXI-Stream Transmit Memory Data

    do_csum                    : out std_logic;                                       --  Enable to do CSUM
    csum_result                : out std_logic_vector(15 downto 0);                   --  Final CSUM result valid with csum_en
    csum_en                    : out std_logic;                                       --  Final CSUM resullt is valid
    csum_we                    : out std_logic_vector(3 downto 0);                    --  Memory Write Enables for 16-bit access
    csum_cmplt                 : out std_logic                                        --  Current CSUM calculation is complete
  );

end tx_csum_partial_calc_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of tx_csum_partial_calc_if is

signal do_csum_int           : std_logic;
signal csum_byte_3_2_en      : std_logic;
signal csum_byte_1_0_en      : std_logic;
signal csum_started          : std_logic;
signal csum_result_int       : std_logic_vector(15 downto 0);

signal csum_3_2              : unsigned(16 downto 0);
signal csum_1_0              : unsigned(16 downto 0);
signal csum_we_int           : std_logic_vector( 3 downto 0);
signal csum_en_int           : std_logic;
signal inc_txd_addr_one_dly1 : std_logic;
signal inc_txd_addr_one_dly2 : std_logic;
signal inc_txd_addr_one_dly3 : std_logic;
signal inc_txd_addr_one_dly4 : std_logic;
signal csum_clr              : std_logic;
signal csum_cmplt_int        : std_logic;

begin

GEN_LEGACY_CSUM : if C_TXCSUM = 1 generate
begin

  CSUM_ENABLE : process(AXI_STR_TXC_ACLK)
  begin

    if rising_edge(AXI_STR_TXC_ACLK) then
      if reset2axi_str_txc = '1' then
        do_csum_int <= '0';
      else
        if axi_str_txc_tready_int_dly = '1' and
           axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tlast_dly0 = '1' then
          case axi_flag is
            when "1010" =>
              case csum_cntrl is
                when "01"   => do_csum_int <= '1';
                when others => do_csum_int <= '0';
              end case;
            when others =>
              do_csum_int <= '0';
          end case;
        else
          do_csum_int <= do_csum_int;
        end if;
      end if;
    end if;
  end process;

  do_csum <= do_csum_int;


-------------------------------------------------------------------------------
--  The legacy CSUM stipulates that the starting position must be 16 bit
--  aligned
-------------------------------------------------------------------------------
SET_CSUM_ENABLES : process(AXI_STR_TXD_ACLK)
begin

  if rising_edge(AXI_STR_TXD_ACLK) then
    if reset2axi_str_txd = '1' or csum_clr = '1' then
      csum_byte_3_2_en <= '0';
      csum_byte_1_0_en <= '0';
      csum_started     <= '0';
    else
      if csum_addr = csum_begin and inc_txd_wr_addr = '1'then
        if csum_begin_bytes(1) = '1' then
          --  Set the enables for the 16 bit csums for 16 bit alignment
          --    Only enable the lower 16 bit csum for the first clock
          csum_byte_3_2_en <= '1';
          csum_byte_1_0_en <= '0';
          csum_started     <= '1';
        else
          --  Otherwise enable both of them
          csum_byte_3_2_en <= '1';
          csum_byte_1_0_en <= '1';
          csum_started     <= '1';
        end if;
      elsif csum_started = '1' and inc_txd_wr_addr = '1' then
        --  once started keep the enables asserted until the end
        --  of the packet
        csum_byte_3_2_en <= '1';
        csum_byte_1_0_en <= '1';
        csum_started     <= '1';
      else
        csum_byte_3_2_en <= csum_byte_3_2_en;
        csum_byte_1_0_en <= csum_byte_1_0_en;
        csum_started     <= csum_started    ;
      end if;
    end if;
  end if;
end process;

DELAY_END_CSUM : process(AXI_STR_TXD_ACLK)
begin

  if rising_edge(AXI_STR_TXD_ACLK) then
    inc_txd_addr_one_dly1 <= inc_txd_addr_one;
    inc_txd_addr_one_dly2 <= inc_txd_addr_one_dly1;
    inc_txd_addr_one_dly3 <= inc_txd_addr_one_dly2;
    inc_txd_addr_one_dly4 <= inc_txd_addr_one_dly3;
    csum_clr              <= inc_txd_addr_one_dly4;
  end if;
end process;




BYTE_3_2_CSUM : process(AXI_STR_TXD_ACLK)
begin

  if rising_edge(AXI_STR_TXD_ACLK) then
    if reset2axi_str_txd = '1' then
      csum_3_2 <= (others => '0');
    else
      if load_csum_int = '1' then
      --  Need to byte swap to properly offset the initial value
        csum_3_2 <= unsigned('0' & csum_init(7 downto 0) & csum_init(15 downto 8));
      elsif inc_txd_addr_one_dly1 = '1' then
      --  add the carry at the end of the csum calculation
         csum_3_2 <= ('0' & csum_3_2(15 downto 0)) + (X"0000" & csum_3_2(16));
      elsif csum_byte_3_2_en = '1' and
            (inc_txd_wr_addr = '1' or inc_txd_addr_one = '1' or non_xilinx_ip_pulse = '1') then
      --  continually calculate the csum for each 16 bits written to memory
        csum_3_2 <= ('0' & csum_3_2(15 downto 0)) +                         -- always zero out the carry
                    unsigned('0' & axi_str_txd_tdata_dly1(31 downto 16)) +  -- add the data to the csum
                    (X"0000" & csum_3_2(16));                               -- add the carry when it occurs
      else
        csum_3_2 <= csum_3_2;
      end if;
    end if;
  end if;
end process;


BYTE_1_0_CSUM : process(AXI_STR_TXD_ACLK)
begin

  if rising_edge(AXI_STR_TXD_ACLK) then
    if reset2axi_str_txd = '1' or csum_clr = '1' then
      csum_1_0 <= (others => '0');
    else
      if inc_txd_addr_one_dly2 = '1' then
      --  Both csum_3_2 and csum_1_0 are calculated, but they need to be added
      --    to each other and then checked for overflow (inc_txd_addr_one_dly2)
         csum_1_0 <= ('0' & csum_3_2(15 downto 0)) + ('0' & csum_1_0(15 downto 0));
      elsif inc_txd_addr_one_dly1 = '1' or inc_txd_addr_one_dly3 = '1' then
      --  add the carry at the end of the data written to memory or
      --  add the carry at the end of the csum calculation
      --    (after csum 3_2 has been added to csum(1_0))
         csum_1_0 <= ('0' & csum_1_0(15 downto 0)) + (X"0000" & csum_1_0(16));
      elsif csum_byte_1_0_en = '1' and
            (inc_txd_wr_addr = '1' or inc_txd_addr_one = '1' or non_xilinx_ip_pulse = '1') then
      --  continually calculate the csum for each 16 bits written to memory
        csum_1_0 <= ('0' & csum_1_0(15 downto 0)) +                          -- always zero out the carry
                    unsigned('0' & axi_str_txd_tdata_dly1(15 downto  0)) +  -- add the data to the csum
                    (X"0000" & csum_1_0(16));                               -- add the carry when it occurs
      else
        csum_1_0 <= csum_1_0;
      end if;
    end if;
  end if;
end process;


--  There is not way of detecting TCP or UDP with legacy CSUM, so always treat it as UDP
--    ie if csum_1_0 = x"FFFF" then invert it.

--  The requirement for checksum is to invert the final value, if it is "0x0000" then
--  set it back to "0xFFFF".  To save a step of inversion, just check it to see if it is
--  0xFFFF before the inversion, and if it is, then do not invert it.

  csum_result_int <= x"FFFF" when (inc_txd_addr_one_dly4 = '1' and csum_1_0 = x"FFFF") else
                     not std_logic_vector(csum_1_0(15 downto 0));

  csum_we_int <= "1100" when inc_txd_addr_one_dly4 = '1' and csum_insert_bytes(1) = '1' else
                 "0011" when inc_txd_addr_one_dly4 = '1' and csum_insert_bytes(1) = '0' else
                 "0000";

  csum_en_int <= '1' when (do_csum_int = '1' and inc_txd_addr_one_dly4 = '1') else
                 '0';


  csum_en     <= csum_en_int;
  csum_we     <= csum_we_int;
  csum_result <= csum_result_int;


  CSUM_COMPLETE : process(AXI_STR_TXD_ACLK)
  begin

    if rising_edge(AXI_STR_TXD_ACLK) then
      if reset2axi_str_txd = '1' then
        csum_cmplt_int <= '0';
      else
        if do_csum_int = '1' then
          if inc_txd_addr_one_dly3 = '1' then
            csum_cmplt_int <= '1';
          else
            csum_cmplt_int <= '0';
          end if;
        else
          if inc_txd_addr_one = '1' then
            csum_cmplt_int <= '1';
          else
            csum_cmplt_int <= '0';
          end if;
        end if;
      end if;
    end if;
  end process;

  csum_cmplt  <= csum_cmplt_int;

end generate GEN_LEGACY_CSUM;



GEN_FULL_CSUM : if C_TXCSUM = 2 generate
begin

  CSUM_ENABLE : process(AXI_STR_TXC_ACLK)
  begin

    if rising_edge(AXI_STR_TXC_ACLK) then
      if reset2axi_str_txc = '1' then
        do_csum_int <= '0';
      else
        if axi_str_txc_tready_int_dly = '1' and
           axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tlast_dly0 = '1' then
          case axi_flag is
            when "1111" =>
              case csum_cntrl is
                when "10"   => do_csum_int <= '1';
                when others => do_csum_int <= '0';
              end case;
            when others =>
              do_csum_int <= '0';
          end case;
        else
          do_csum_int <= do_csum_int;
        end if;
      end if;
    end if;
  end process;

do_csum     <= '0';
csum_result <= (others => '0');
csum_en     <= '0';
csum_we     <= (others => '0');
csum_cmplt  <= '1';

end generate GEN_FULL_CSUM;


end rtl;


-------------------------------------------------------------------------------
-- tx_csum_full_fsm - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_csum_full_fsm.vhd
-- Version:         v1.00a
-- Description:     top level of embedded ip Ethernet MAC interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--                    tx_axistream_if.vhd
--                      tx_basic_if.vhd
--                      tx_csum_if.vhd
--                        tx_csum_full_if.vhd
--          ->              tx_csum_full_fsm.vhd
--                          tx_csum_full_calc_if.vhd
--                        tx_partial_csum_if.vhd
--                          tx_csum_partial_calc_if.vhd
--                      tx_vlan_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tx_if_pack.all;



-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity tx_csum_full_fsm is
  generic (
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32     := 32;
    c_TxD_addrb_width      : integer range  0 to 13     := 10
  );
  port (

    AXI_STR_TXD_ACLK  : in  std_logic;                                        --  Clock
    reset2axi_str_txd : in  std_logic;                                        --  Reset

    txd_strbs         : in  std_logic_vector(3 downto 0);                     --  AXI-Stream Tx Data Strobes
    do_csum           : in  std_logic;                                        --  axi_flag must = 0xA for this to be enabled
    abort_csum        : out std_logic;                                        --  All conditions were not met to complete csum
    txd_tlast         : in  std_logic;                                        --  AXI-Stream Tx Data Last
    csum_calc_en      : in  std_logic;                                        --  axi_str_txd_tvalid_dly0 and
                                                                              --  axi_str_txd_tready_int_dly;
    clr_csums         : out std_logic;                                        --  Clear CSUM flags and calculations
    tcp_ptcl          : out std_logic;                                        --  TCP Protocol Indicator
    udp_ptcl          : out std_logic;                                        --  UDP Protocol Indicator
    en_ipv4_hdr_b32   : out std_logic_vector( 1 downto 0);                    --  bytes 3 and 2 of din
    en_ipv4_hdr_b10   : out std_logic_vector( 1 downto 0);                    --  bytes 1 and 0 of din
    last_ipv4_hdr_cnt : out std_logic;                                        --  last data for IPv4 Header Calculation
    fsm_csum_en_b32   : out std_logic_vector( 1 downto 0);                    --  bytes 3 and 2 of din
    fsm_csum_en_b10   : out std_logic_vector( 1 downto 0);                    --  bytes 1 and 0 of din
    add_psdo_wd       : out std_logic;                                        --  last data for TCP/UDP Calculation
    ptcl_csum_cmplt   : in  std_logic;                                        --  indicates the TCP/UDP csum calculation is complete
    zeroes_en         : out std_logic_vector( 1 downto 0);                    --  stalls the CSUM calculations for one clock so
                                                                              --  Zeroes do not need muxed in
    din               : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1  downto 0); --  AXI Stream Tx Data
    csum_din          : out std_logic_vector(C_S_AXI_DATA_WIDTH-1  downto 0); --  Mux out of pseudo data or axi_str_txd_tdata_dly0
    do_ipv4hdr        : out std_logic;                                        --  only do the ipv4 header csum
    not_tcp_udp       : out std_logic;                                        --  only do the ipv4 header csum - no TCP/UDP protocol
    do_full_csum      : out std_logic;                                        --  do the ipv4 headr and TCP/UDP csum
    hdr_csum_cmplt    : in  std_logic;                                        --  Header CSUM Calculation is complete
    wr_hdr_csum       : out std_logic;                                        --  Enable to Write the Header CSUM to Memory
    wr_ptcl_csum      : out std_logic;                                        --  Enable to Write the EthII/Snap Ipv4 TCP/UDP CSUM

    csum_strt_addr    : in  std_logic_vector(c_TxD_addrb_width-1   downto 0); --  Start Address to start the CSUM ccalculation
    csum_ipv4_hdr_addr: out std_logic_vector(c_TxD_addrb_width-1   downto 0); --  IPv4 Header Start Address
    csum_ipv4_hdr_we  : out std_logic_vector( 3 downto 0);                    --  IPv4 Header Write Enable to Memory
    csum_ptcl_addr    : out std_logic_vector(c_TxD_addrb_width-1   downto 0); --  Address to Write the EthII/Snap Ipv4 TCP/UDP CSUM
    csum_ptcl_we      : out std_logic_vector( 3 downto 0)                     --  Enables to Write the EthII/Snap Ipv4 TCP/UDP CSUM


  );

end tx_csum_full_fsm;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of tx_csum_full_fsm is

  signal din_big_end           : std_logic_vector(0 to C_S_AXI_DATA_WIDTH-1);

  type   FULL_CSUM_FSM_TYPE is (
           IDLE,
           DST,     --  Destination Address
           DST_SRC, --  Destination and Source Address
           SRC,     --  Source Address
           IDF,     --  Identify Frame Type
           SNAP,    --  SNAP Frame
           OUI,     --  SNAP OUI
           IPV4_HDR,--  IPv4 Header
           PCOL_HDR,--  Protocol of the packet - TCP or UDP
           DATA,    --  Data
           WAIT_TLAST,
           WR_HDR_ONLY,
           WAIT_DELAY,
           WAIT_COMPLETE,
           WR_HDR,  --  Write Header CSUM
           WR_CSUM  --  Write TCP/UDP CSUM
           );
  signal fcsum_wr_cs, fcsum_wr_ns             : FULL_CSUM_FSM_TYPE;

  signal store_hdr_length     : std_logic;
  signal hdr_length           : unsigned( 5 downto 0);

  signal en_ipv4_hdr_cnt      : std_logic;
  signal en_ipv4_hdr_b10_int  : std_logic_vector(1 downto 0);
  signal en_ipv4_hdr_b32_int  : std_logic_vector(1 downto 0);



  signal clr_hdr_cnt          : std_logic;
  signal last_ipv4_hdr_cnt_int: std_logic;
  signal en_pcol_hdr_cnt      : std_logic;
  signal hdr_cnt              : unsigned( 2 downto 0);
  signal store_version        : std_logic;
  signal version              : std_logic_vector( 3 downto 0);
  signal calc_frm_length      : std_logic;
  signal frm_length           : std_logic_vector(0 to 15);
  signal fsm_csum_en          : std_logic;
  signal fsm_csum_en_b32_int  : std_logic_vector(1 downto 0);
  signal fsm_csum_en_b10_int  : std_logic_vector(1 downto 0);

  signal csum_ipv4_hdr_addr_int : unsigned(c_TxD_addrb_width-1   downto 0);
  signal csum_ipv4_hdr_we_int : std_logic_vector( 3 downto 0);
  signal csum_ptcl_addr_int   : unsigned(c_TxD_addrb_width-1   downto 0);
  signal csum_ptcl_we_int     : std_logic_vector( 3 downto 0);

  signal store_sa_da          : std_logic;
  signal sa0                  : std_logic_vector(15 downto 0); --Source Address Half word - Little End
  signal sa1                  : std_logic_vector(15 downto 0); --Source Address Half word - Little End
  signal da0                  : std_logic_vector(15 downto 0); --Destination Address Half word - Little End
  signal da1                  : std_logic_vector(15 downto 0); --Destination Address Half word - Little End
  signal clr_csums_int        : std_logic;



  signal set_eth2             : std_logic;
  signal eth2                 : std_logic;
  signal set_snap             : std_logic;
  signal snap_hit             : std_logic;
  signal set_oui_hit          : std_logic;
  signal oui_hit              : std_logic;
  signal set_vlan             : std_logic;
  signal vlan                 : std_logic;
  signal set_ipv4             : std_logic;
  signal ipv4                 : std_logic;
  signal set_ptcl             : std_logic;
  signal tcp_ptcl_int         : std_logic;
  signal udp_ptcl_int         : std_logic;
  signal set_ipv4hdr_only     : std_logic;
  signal do_ipv4_int          : std_logic;

  signal set_fragment         : std_logic;
  signal fragment             : std_logic;

  signal do_full_csum_int     : std_logic;
  signal add_psdo_wd_int      : std_logic;
  signal pseudo_data          : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal zeroes_en_int        : std_logic_vector(1 downto 0);

  signal abort_csum_int       : std_logic;

  signal set_not_tcp_udp      : std_logic;
  signal not_tcp_udp_int      : std_logic;

  begin

    clr_csums           <= clr_csums_int;
    tcp_ptcl            <= tcp_ptcl_int;
    udp_ptcl            <= udp_ptcl_int;
    do_ipv4hdr          <= do_ipv4_int;
    not_tcp_udp         <= not_tcp_udp_int;
    do_full_csum        <= do_full_csum_int;

    en_ipv4_hdr_b32     <= en_ipv4_hdr_b32_int;
    en_ipv4_hdr_b10     <= en_ipv4_hdr_b10_int;
    last_ipv4_hdr_cnt   <= last_ipv4_hdr_cnt_int;
    fsm_csum_en_b32     <= fsm_csum_en_b32_int;
    fsm_csum_en_b10     <= fsm_csum_en_b10_int;
    add_psdo_wd         <= add_psdo_wd_int;
    zeroes_en           <= zeroes_en_int;

    csum_ipv4_hdr_addr  <= std_logic_vector(csum_ipv4_hdr_addr_int);
    csum_ipv4_hdr_we    <= csum_ipv4_hdr_we_int;
    csum_ptcl_addr      <= std_logic_vector(csum_ptcl_addr_int);
    csum_ptcl_we        <= csum_ptcl_we_int;

    -- Little endian to Big Endian
    din_big_end( 0 to  7) <= din( 7 downto  0);
    din_big_end( 8 to 15) <= din(15 downto  8);
    din_big_end(16 to 23) <= din(23 downto 16);
    din_big_end(24 to 31) <= din(31 downto 24);



    -----------------------------------------------------------------------
    --  FSM used to control the Full Checksum calculation
    -----------------------------------------------------------------------
    FSM_FULL_CSUM_CMB : process(fcsum_wr_cs,csum_calc_en,do_csum,
      din,din_big_end,
      vlan,hdr_cnt,ipv4,eth2,snap_hit,oui_hit,
      udp_ptcl_int,tcp_ptcl_int,fragment,
      txd_tlast,ptcl_csum_cmplt,txd_strbs,hdr_csum_cmplt,
      not_tcp_udp_int,do_ipv4_int
      )

    begin

      store_hdr_length     <= '0';
      en_ipv4_hdr_cnt      <= '0';
      en_ipv4_hdr_b10_int  <= "00";
      en_ipv4_hdr_b32_int  <= "00";

      last_ipv4_hdr_cnt_int<= '0';
      en_pcol_hdr_cnt      <= '0';
      clr_hdr_cnt          <= '0';
      store_version        <= '0';
      calc_frm_length      <= '0';
      fsm_csum_en          <= '0';
      fsm_csum_en_b32_int  <= "00";
      fsm_csum_en_b10_int  <= "00";

      store_sa_da          <= '0';
      wr_hdr_csum          <= '0';
      wr_ptcl_csum         <= '0';
      clr_csums_int        <= '0';

      set_eth2             <= '0';
      set_snap             <= '0';
      set_oui_hit          <= '0';
      set_vlan             <= '0';
      set_ipv4             <= '0';
      set_ptcl             <= '0';
      set_ipv4hdr_only     <= '0';

      set_fragment         <= '0';
      zeroes_en_int        <= "00";

      add_psdo_wd_int      <= '0';

      abort_csum_int       <= '0';

      set_not_tcp_udp      <= '0';

      case fcsum_wr_cs is
        when IDLE      =>
          if do_csum = '1' and csum_calc_en = '1' then
          --  Flag is set and tvalid/tready are HIGH
          --  If csum calc is aborted because all conditions are not met
          --    (not IPv4, not TCP, not UDP, etc) then do_csum is cleared
          --    which will prevent the FSM from starting again until the next packet
            fcsum_wr_ns <= DST;
          else
            fcsum_wr_ns <= IDLE;
          end if;
        when DST      =>
          if csum_calc_en = '1' then
          --  tvalid/tready are HIGH
            fcsum_wr_ns <= DST_SRC;
          else
            fcsum_wr_ns <= DST;
          end if;
        when DST_SRC  =>
          if csum_calc_en = '1' then
          --  tvalid/tready are HIGH
            fcsum_wr_ns <= SRC;
          else
            fcsum_wr_ns <= DST_SRC;
          end if;
        when SRC      =>
          if txd_tlast = '1' and csum_calc_en = '1' then
            --  Tlast was received so exit
            clr_csums_int       <= '0';
            abort_csum_int      <= '0';
            add_psdo_wd_int     <= '1';         --  pseudo word is not done, but this needs to set
                                                --  ptcl_csum_cmplt and exit tx_csum_full_if.vhd FSMs
            fcsum_wr_ns         <= WAIT_COMPLETE;
          elsif csum_calc_en = '1' then
            if din(15 downto 0) = X"0081" then
            --  It is VLAN
              set_vlan         <= '1';
              set_snap         <= '0';
              set_eth2         <= '0';
              store_hdr_length <= '0';
              en_ipv4_hdr_cnt  <= '0';
              store_version    <= '0';
              set_ipv4         <= '0';
              fcsum_wr_ns      <= IDF;
            elsif din_big_end(0 to 15) <= X"0600" and   --Length is less than 0x600 and
                  din(23 downto 16)  = X"AA" and din(31 downto 24) = X"AA"  then --DSAP and SSAP
            --  It is SNAP
              set_vlan         <= '0';
              set_snap         <= '1';
              set_eth2         <= '0';
              store_hdr_length <= '0';
              en_ipv4_hdr_cnt  <= '0';
              store_version    <= '0';
              set_ipv4         <= '0';
              fcsum_wr_ns      <= IDF;  --
            elsif din(15 downto  0) = X"0008" and -- TYPE is 0x0800 (IPv4) and
                  din(23 downto 16) = X"45" then  -- Version = 0x4 (IPv4) and HDR Length = 5
            -- It is Ethernet II IPv4 with 5 word header  -- IPv4 header options are not supported
              set_vlan             <= '0';
              set_snap             <= '0';
              set_eth2             <= '1';
              store_hdr_length     <= '1';  --  length of packet starting from here, to the end (+4 words for EII, +1+ vlan, +2 snap
              en_ipv4_hdr_cnt      <= '1';
              en_ipv4_hdr_b10_int  <= "00";
              en_ipv4_hdr_b32_int  <= "11";
              store_version        <= '1';
              set_ipv4             <= '1';
              fcsum_wr_ns          <= IPV4_HDR;


            else -- Not all conditions were met to perform CSUM
              set_vlan             <= '0';
              set_snap             <= '0';
              set_eth2             <= '0';
              store_hdr_length     <= '0';
              en_ipv4_hdr_cnt      <= '0';
              en_ipv4_hdr_b10_int  <= "00";
              en_ipv4_hdr_b32_int  <= "00";
              store_version        <= '0';
              set_ipv4             <= '0';
              clr_csums_int        <= '0';
              abort_csum_int       <= '0';
              fcsum_wr_ns          <= WAIT_TLAST;--WAIT_COMPLETE;
            end if;
          else
            set_vlan             <= '0';
            set_snap             <= '0';
            set_eth2             <= '0';
            store_hdr_length     <= '0';
            en_ipv4_hdr_cnt      <= '0';
            en_ipv4_hdr_b10_int  <= "00";
            en_ipv4_hdr_b32_int  <= "00";
            store_version        <= '0';
            set_ipv4             <= '0';
            fcsum_wr_ns          <= SRC;
          end if;
        when IDF =>
          if txd_tlast = '1' and csum_calc_en = '1' then
            --  Tlast was received so exit
            clr_csums_int       <= '0';
            abort_csum_int      <= '0';
            add_psdo_wd_int     <= '1';         --  pseudo word is not done, but this needs to set
                                                --  ptcl_csum_cmplt and exit tx_csum_full_if.vhd FSMs
            fcsum_wr_ns         <= WAIT_COMPLETE;
          elsif csum_calc_en = '1' then
            if vlan = '1' then
              if din(15 downto 0) = X"0008" and  -- TYPE is 0x0800 (IPv4) and
                 din(23 downto 16) = X"45" then  -- Version = 0x4 (IPv4) and HDR Length = 5
                -- It is Ethernet II IPv4 with 5 word header
                store_hdr_length     <= '1';
                en_ipv4_hdr_cnt      <= '1';
                en_ipv4_hdr_b10_int  <= "00";
                en_ipv4_hdr_b32_int  <= "11";
                store_version        <= '1';
                set_eth2             <= '1';
                set_ipv4             <= '1';
                set_snap             <= '0';
                fcsum_wr_ns          <= IPV4_HDR;
              elsif din_big_end(0 to 15) <= X"0600" and  -- Length is less than 0x600 and
                  din(23 downto 16) = X"AA" and din(31 downto 24) = X"AA" then --DSAP and SSAP
                -- It is Ethernet SNAP
                store_hdr_length <= '0';
                en_ipv4_hdr_cnt  <= '0';
                store_version    <= '0';
                set_eth2         <= '0';
                set_ipv4         <= '0';
                set_snap         <= '1';
                fcsum_wr_ns      <= SNAP;  -- SNAP detected so check OUI
              else
                store_hdr_length <= '0';
                en_ipv4_hdr_cnt  <= '0';
                store_version    <= '0';
                set_eth2         <= '0';
                set_ipv4         <= '0';
                set_snap         <= '0';
                clr_csums_int    <= '0';
                abort_csum_int   <= '0';
                fcsum_wr_ns      <= WAIT_TLAST;--WAIT_COMPLETE;  -- Do not do CSUM
              end if;
            else -- eth_snap_xsap_hit = '1' then
              if din( 7 downto  0) = X"03" and  -- Endian Swap  -- Control
                 din(15 downto  8) = X"00" and  -- Endian Swap  -- OUI
                 din(23 downto 16) = X"00" and  -- Endian Swap  -- OUI
                 din(31 downto 24) = X"00" then -- Endian Swap  -- OUI
                store_hdr_length <= '0';
                en_ipv4_hdr_cnt  <= '0';
                store_version    <= '0';
                set_eth2         <= '0';
                set_ipv4         <= '0';
                set_snap         <= '0';
                set_oui_hit      <= '1';
                fcsum_wr_ns      <= OUI;
              else
                store_hdr_length <= '0';
                en_ipv4_hdr_cnt  <= '0';
                store_version    <= '0';
                set_eth2         <= '0';
                set_ipv4         <= '0';
                set_snap         <= '0';
                set_oui_hit      <= '0';
                clr_csums_int    <= '0';
                abort_csum_int   <= '0';
                fcsum_wr_ns      <= WAIT_TLAST;--WAIT_COMPLETE;
              end if;
            end if;
          else
            set_eth2         <= '0';
            set_ipv4         <= '0';
            set_snap         <= '0';
            set_oui_hit      <= '0';
            fcsum_wr_ns      <= IDF;
          end if;
        when SNAP =>
          if txd_tlast = '1' and csum_calc_en = '1' then
            --  Tlast was received so exit
            clr_csums_int       <= '0';
            abort_csum_int      <= '0';
            add_psdo_wd_int     <= '1';         --  pseudo word is not done, but this needs to set
                                                --  ptcl_csum_cmplt and exit tx_csum_full_if.vhd FSMs
            fcsum_wr_ns         <= WAIT_COMPLETE;
          elsif csum_calc_en = '1' then
            if din( 7 downto  0) = X"03" and  -- Control
               din(15 downto  8) = X"00" and  -- OUI
               din(23 downto 16) = X"00" and  -- OUI
               din(31 downto 24) = X"00" then -- OUI
              set_oui_hit      <= '1';
              fcsum_wr_ns      <= OUI;
            else --was not OUI hit or last was received so exit
              set_oui_hit      <= '0';
              clr_csums_int    <= '0';
              abort_csum_int   <= '0';
              fcsum_wr_ns      <= WAIT_TLAST;--WAIT_COMPLETE;
            end if;
          else
            set_oui_hit      <= '0';
            fcsum_wr_ns      <= SNAP;
          end if;
        when OUI =>
          if txd_tlast = '1' and csum_calc_en = '1' then
            --  Tlast was received so exit
            clr_csums_int       <= '0';
            abort_csum_int      <= '0';
            add_psdo_wd_int     <= '1';         --  pseudo word is not done, but this needs to set
                                                --  ptcl_csum_cmplt and exit tx_csum_full_if.vhd FSMs
            fcsum_wr_ns         <= WAIT_COMPLETE;
          elsif csum_calc_en = '1' then

            if din(15 downto 0) = X"0008" and  -- TYPE is 0x0800 (IPv4) and
               din(23 downto 16) = X"45" then    -- It is SNAP IPv4 with 5 word header
              store_hdr_length     <= '1';
              en_ipv4_hdr_cnt      <= '1';
              en_ipv4_hdr_b10_int  <= "00";
              en_ipv4_hdr_b32_int  <= "11";
              store_version        <= '1';
              set_ipv4             <= '1';
              clr_csums_int        <= '0';
              abort_csum_int       <= '0';
              fcsum_wr_ns          <= IPV4_HDR;
            else --  Not ipv4 so go to idle
              store_hdr_length     <= '0';
              en_ipv4_hdr_cnt      <= '0';
              en_ipv4_hdr_b10_int  <= "00";
              en_ipv4_hdr_b32_int  <= "00";
              store_version        <= '0';
              set_ipv4             <= '0';
              clr_csums_int        <= '0';
              abort_csum_int       <= '0';
              fcsum_wr_ns          <= WAIT_TLAST;--WAIT_COMPLETE;
            end if;

          else
            store_hdr_length     <= '0';
            en_ipv4_hdr_cnt      <= '0';
            en_ipv4_hdr_b10_int  <= "00";
            en_ipv4_hdr_b32_int  <= "00";
            store_version        <= '0';
            set_ipv4             <= '0';
            clr_csums_int        <= '0';
            abort_csum_int       <= '0';
            fcsum_wr_ns          <= OUI;
          end if;
        when IPV4_HDR =>
          if csum_calc_en = '1' then
            case hdr_cnt is
              when "001" => calc_frm_length     <= '1';
                            set_ptcl            <= '0';
                            store_sa_da         <= '0';
                            fsm_csum_en         <= '0';
                            en_ipv4_hdr_cnt     <= '1';
                            en_ipv4_hdr_b10_int <= "11";
                            en_ipv4_hdr_b32_int <= "11";
                            clr_hdr_cnt         <= '0';
                            fcsum_wr_ns         <= IPV4_HDR;
              when "010" => calc_frm_length     <= '0';
                            set_ptcl            <= '1';
                            store_sa_da         <= '0';
                            fsm_csum_en         <= '0';
                            en_ipv4_hdr_cnt     <= '1';
                            en_ipv4_hdr_b10_int <= "11";
                            en_ipv4_hdr_b32_int <= "11";
                            clr_hdr_cnt         <= '0';
                            fcsum_wr_ns         <= IPV4_HDR;
                            if --din(6) = '1' and --  Don't Fragment (DF) = '1'
                               din(5) = '0' and --  More Fragment (MF) Flag = '0'
                               din(4) = '0' and               -- Fragment Offset
                               din(3 downto 0) = X"0" and     -- Fragment Offset
                               din(15 downto  8) = X"00" then -- Fragment Offset
                              set_fragment <= '0';
                            else
                              set_fragment <= '1';
                            end if;
              when "011" => --  mw 1220 --  if ipv4 = '1' and
                            --  mw 1220 --     (eth2 = '1' or (snap_hit = '1' and oui_hit = '1')) then --and
                -- two types of ipv4 frames Ethernet II and SNAP
                            --  Check to ensure all conditions are met before
                            --  continuing with csum
                              calc_frm_length     <= '0';
                              set_ptcl            <= '0';
                              store_sa_da         <= '1';
                              fsm_csum_en         <= '1';
                              fsm_csum_en_b32_int <= "11";
                              fsm_csum_en_b10_int <= "00";
                              en_ipv4_hdr_cnt     <= '1';
                              en_ipv4_hdr_b10_int <= "11";
                              en_ipv4_hdr_b32_int <= "11";
                              zeroes_en_int       <= "01";  -- Set enable for ipv4 header csum to insert zeroes into calculation
                              clr_hdr_cnt         <= '0';
                              clr_csums_int       <= '0';
                              abort_csum_int      <= '0';
                              fcsum_wr_ns         <= IPV4_HDR;
             when "100" =>  calc_frm_length       <= '0';
                            set_ptcl              <= '0';
                            store_sa_da           <= '1';
                            fsm_csum_en           <= '1';
                            fsm_csum_en_b32_int   <= "11";
                            fsm_csum_en_b10_int   <= "11";
                            en_ipv4_hdr_cnt       <= '1';
                            en_ipv4_hdr_b10_int   <= "11";
                            en_ipv4_hdr_b32_int   <= "11";
                            last_ipv4_hdr_cnt_int <= '0';
                            clr_hdr_cnt           <= '1';
                            if (tcp_ptcl_int = '1' or udp_ptcl_int = '1') and fragment = '0' then
                              set_ipv4hdr_only <= '0';
                              set_not_tcp_udp  <= '0';
                              fcsum_wr_ns      <= PCOL_HDR;
                            else -- Only perform the IPv4 Header CSUM -- Only IPv4 is set
                              set_ipv4hdr_only <= '1';
                              set_not_tcp_udp  <= '1';
                              fcsum_wr_ns      <= WAIT_TLAST;--WR_HDR_ONLY;
                           end if;
              when others=> calc_frm_length       <= '0';
                            set_ptcl              <= '0';
                            store_sa_da           <= '0';
                            fsm_csum_en           <= '0';
                            fsm_csum_en_b32_int   <= "00";
                            fsm_csum_en_b10_int   <= "00";
                            en_ipv4_hdr_cnt       <= '0';
                            en_ipv4_hdr_b10_int   <= "00";
                            en_ipv4_hdr_b32_int   <= "00";
                            clr_hdr_cnt           <= '0';
                            fcsum_wr_ns           <= IPV4_HDR;
            end case;
          else
            calc_frm_length     <= '0';
            set_ptcl            <= '0';
            store_sa_da         <= '0';
            fsm_csum_en         <= '0';
            fsm_csum_en_b32_int <= "00";
            fsm_csum_en_b10_int <= "00";
            en_ipv4_hdr_cnt     <= '0';
            en_ipv4_hdr_b10_int <= "00";
            en_ipv4_hdr_b32_int <= "00";
            clr_hdr_cnt         <= '0';
            fcsum_wr_ns         <= IPV4_HDR;
          end if;
        when PCOL_HDR =>

          if csum_calc_en = '1' then
            fsm_csum_en         <= '1';
            fsm_csum_en_b32_int <= "11";
            fsm_csum_en_b10_int <= "11";
            case hdr_cnt is
            --  when TCP this count will reset after "100"
            --  when udp this count will reset after "001"
              when "000" => calc_frm_length       <= '0';
                            store_sa_da           <= '1';
                            en_ipv4_hdr_cnt       <= '0';
                            en_ipv4_hdr_b10_int   <= "11";
                            en_ipv4_hdr_b32_int   <= "00";
                            last_ipv4_hdr_cnt_int <= '1';
                            en_pcol_hdr_cnt       <= '1';
                            zeroes_en_int         <= "00";
                            fcsum_wr_ns           <= PCOL_HDR;
              when "001" => if udp_ptcl_int = '1' then --and fragment = '0' then
                              en_pcol_hdr_cnt <= '0';
                              clr_hdr_cnt     <= '1';
                              calc_frm_length <= '1';
                              zeroes_en_int   <= "00";
                              fcsum_wr_ns     <= DATA;
                            elsif tcp_ptcl_int = '1' then --and fragment = '0' then --has to be TCP
                              en_pcol_hdr_cnt <= '1';
                              clr_hdr_cnt     <= '0';
                              calc_frm_length <= '0';
                              zeroes_en_int   <= "00";
                              fcsum_wr_ns     <= PCOL_HDR;
                            else -- it was not IPv4, tcp/udp, and fragments /= 0
                              en_pcol_hdr_cnt <= '0';
                              clr_hdr_cnt     <= '0';
                              zeroes_en_int   <= "00";
                              clr_csums_int   <= '0';
                              abort_csum_int  <= '0';
                              fcsum_wr_ns     <= WAIT_TLAST;--WAIT_COMPLETE;
                            end if;
              when "100" => en_pcol_hdr_cnt <= '0';
                            clr_hdr_cnt     <= '1';
                            zeroes_en_int   <= "10";  -- Set enable for data csum to insert zeroes into calculation
                            fcsum_wr_ns     <= DATA;

              when others=> en_pcol_hdr_cnt <= '1';
                            clr_hdr_cnt     <= '0';
                            zeroes_en_int   <= "00";
                            fcsum_wr_ns     <= PCOL_HDR;
            end case;
          else
            en_pcol_hdr_cnt     <= '0';
            clr_hdr_cnt         <= '0';
            zeroes_en_int       <= "00";
            fsm_csum_en         <= '0';
            fsm_csum_en_b32_int <= "00";
            fsm_csum_en_b10_int <= "00";
            fcsum_wr_ns         <= PCOL_HDR;
          end if;

        when DATA     =>
          if csum_calc_en = '1' and udp_ptcl_int = '1' and hdr_cnt = "000" then
            zeroes_en_int   <= "01";
            en_pcol_hdr_cnt <= '1';
          else
            zeroes_en_int   <= "00";
            en_pcol_hdr_cnt <= '0';
          end if;

          if txd_tlast = '1' and csum_calc_en = '1' then
            fsm_csum_en         <= '1';
            fsm_csum_en_b32_int <= txd_strbs(3 downto 2);
            fsm_csum_en_b10_int <= txd_strbs(1 downto 0);
            fcsum_wr_ns         <= WR_HDR;
          elsif txd_tlast = '0' and csum_calc_en = '1' then
            fsm_csum_en         <= '1';
            fsm_csum_en_b32_int <= "11";
            fsm_csum_en_b10_int <= "11";
            fcsum_wr_ns         <= DATA;
          else
            fsm_csum_en         <= '0';
            fsm_csum_en_b32_int <= "00";
            fsm_csum_en_b10_int <= "00";
            fcsum_wr_ns         <= DATA;
          end if;

        when WAIT_TLAST =>
          --  Need to wait for TLAST before completing the CSUM
          if csum_calc_en = '1' then
            case hdr_cnt is
              --  need to assert the header csum enable to include the last bytes
              when "000" =>
                calc_frm_length       <= '0';
                store_sa_da           <= '1';
                en_ipv4_hdr_cnt       <= '0';
                en_ipv4_hdr_b10_int   <= "11";
                en_ipv4_hdr_b32_int   <= "00";
                last_ipv4_hdr_cnt_int <= '1';
                en_pcol_hdr_cnt       <= '1';
                zeroes_en_int         <= "00";
                clr_hdr_cnt           <= '0';
                clr_csums_int         <= '0';
                abort_csum_int        <= '0';
              when others =>
                calc_frm_length       <= '0';
                store_sa_da           <= '0';
                en_ipv4_hdr_cnt       <= '0';
                en_ipv4_hdr_b10_int   <= "00";
                en_ipv4_hdr_b32_int   <= "00";
                last_ipv4_hdr_cnt_int <= '0';
                en_pcol_hdr_cnt       <= '0';
                zeroes_en_int         <= "00";
                clr_hdr_cnt           <= '0';
                clr_csums_int         <= '0';
                abort_csum_int        <= '0';
            end case;
          else
            calc_frm_length       <= '0';
            store_sa_da           <= '0';
            en_ipv4_hdr_cnt       <= '0';
            en_ipv4_hdr_b10_int   <= "00";
            en_ipv4_hdr_b32_int   <= "00";
            last_ipv4_hdr_cnt_int <= '0';
            en_pcol_hdr_cnt       <= '0';
            zeroes_en_int         <= "00";
            clr_hdr_cnt           <= '0';
            clr_csums_int         <= '0';
            abort_csum_int        <= '0';
          end if;

          if txd_tlast = '1' and csum_calc_en = '1' then
          --  Do one of two branches depending upon if the ipv4 header csum was calculated or not
            if do_ipv4_int = '1' then
              add_psdo_wd_int     <= '0';
              fcsum_wr_ns         <= WAIT_DELAY;
            else
              add_psdo_wd_int     <= '1';         --  pseudo word is not done, but this needs to set
                                                  --  ptcl_csum_cmplt and exit tx_csum_full_if.vhd FSMs
              fcsum_wr_ns         <= WAIT_COMPLETE;
            end if;
          else
            fcsum_wr_ns         <= WAIT_TLAST;
          end if;

        when WAIT_DELAY =>
        --  need to delay 1 clock so inc_txd_wr_one does not occur with wr_hdr_csum
          fcsum_wr_ns         <= WR_HDR_ONLY;

        when WR_HDR_ONLY =>
--          --  Got here from IPV4_HDR state so need to enable en_ipv4_hdr_b10_int for last IPv4 header data
--          case hdr_cnt is
--            when "000" =>
--              calc_frm_length       <= '0';
--              store_sa_da           <= '1';
--              en_ipv4_hdr_cnt       <= '0';
--              en_ipv4_hdr_b10_int   <= "11";
--              en_ipv4_hdr_b32_int   <= "00";
--              last_ipv4_hdr_cnt_int <= '1';
--              en_pcol_hdr_cnt       <= '1';
--              zeroes_en_int         <= "00";
--              clr_hdr_cnt           <= '0';
--              clr_csums_int         <= '0';
--              abort_csum_int        <= '0';
--            when others =>
--              calc_frm_length       <= '0';
--              store_sa_da           <= '0';
--              en_ipv4_hdr_cnt       <= '0';
--              en_ipv4_hdr_b10_int   <= "00";
--              en_ipv4_hdr_b32_int   <= "00";
--              last_ipv4_hdr_cnt_int <= '0';
--              en_pcol_hdr_cnt       <= '0';
--              zeroes_en_int         <= "00";
--              clr_hdr_cnt           <= '0';
--              clr_csums_int         <= '0';
--              abort_csum_int        <= '0';
--          end case;

          if hdr_csum_cmplt = '1' then
            wr_hdr_csum         <= '1';
            clr_hdr_cnt         <= '0';
            clr_csums_int       <= '0';
            add_psdo_wd_int     <= '1';           --  pseudo word is not done, but this needs to set
                                                  --  ptcl_csum_cmplt and exit tx_csum_full_if.vhd FSMs
            fcsum_wr_ns         <= WAIT_COMPLETE;
          else
            wr_hdr_csum         <= '0';
            clr_hdr_cnt         <= '0';
            add_psdo_wd_int     <= '0';
            clr_csums_int       <= '0';
            fcsum_wr_ns         <= WR_HDR_ONLY;
          end if;

        when WAIT_COMPLETE   =>
--          if ipv4 = '1' and hdr_cnt = "000" then
--          --  true if got here from IPV4_HDR state
--          --    so enable en_ipv4_hdr_b10_int to get last IPv4 header data
--            calc_frm_length       <= '0';
--            store_sa_da           <= '1';
--            en_ipv4_hdr_cnt       <= '0';
--            en_ipv4_hdr_b10_int   <= "11";
--            en_ipv4_hdr_b32_int   <= "00";
--            last_ipv4_hdr_cnt_int <= '1';
--            en_pcol_hdr_cnt       <= '1';
--            zeroes_en_int         <= "00";
--            clr_hdr_cnt           <= '0';
--            clr_csums_int         <= '0';
--            abort_csum_int        <= '0';
--            fcsum_wr_ns           <= WAIT_COMPLETE;
--          elsif ptcl_csum_cmplt = '1' then
          if ptcl_csum_cmplt = '1' then
            clr_hdr_cnt   <= '1';
            clr_csums_int <= '1';
            abort_csum_int<= '1';
            fcsum_wr_ns   <= IDLE;
          else
            clr_hdr_cnt   <= '0';
            clr_csums_int <= '0';
            abort_csum_int<= '0';
            fcsum_wr_ns   <= WAIT_COMPLETE;
          end if;
        when WR_HDR   =>
          if hdr_csum_cmplt = '1' and (tcp_ptcl_int = '1' or udp_ptcl_int = '1') and fragment = '0' then
            wr_hdr_csum         <= '1';
            clr_csums_int       <= '0';
            add_psdo_wd_int     <= '1';
            fsm_csum_en         <= '1';
            fsm_csum_en_b32_int <= "11";
            fsm_csum_en_b10_int <= "11";
            fcsum_wr_ns         <= WR_CSUM;
          else
            wr_hdr_csum         <= '0';
            clr_csums_int       <= '0';
            add_psdo_wd_int     <= '0';
            fsm_csum_en         <= '0';
            fsm_csum_en_b32_int <= "00";
            fsm_csum_en_b10_int <= "00";
            fcsum_wr_ns         <= WR_HDR;
          end if;
        when WR_CSUM  =>
          if ptcl_csum_cmplt = '1' then
            clr_hdr_cnt  <= '1';
            wr_ptcl_csum <= '1';
            clr_csums_int<= '1';
            fcsum_wr_ns  <= IDLE;
          else
            clr_hdr_cnt  <= '0';
            wr_ptcl_csum <= '0';
            clr_csums_int<= '0';
            fcsum_wr_ns  <= WR_CSUM;
          end if;
        when others =>
          fcsum_wr_ns  <= IDLE;
      end case;
    end process;

    -----------------------------------------------------------------------
    --  FSM Sequencer
    -----------------------------------------------------------------------
    FSM_FULL_CSUM_SEQ : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          fcsum_wr_cs <= IDLE;
        else
          fcsum_wr_cs <= fcsum_wr_ns;
        end if;
      end if;
    end process;



    ---------------------------------------------------------------------------
    --  At store_hdr_length, din contains the header length in words...
    --  Convert it to bytes
    --    IPv4 Header options are not currently supported, so this must
    --    equal 0x5wds (0x14bytes) for the CSUM to be calculated
    ---------------------------------------------------------------------------
    ETHERNET_HEADER_LENGTH_REG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          hdr_length <= (others => '0');
        else
          if store_hdr_length = '1' then
            hdr_length <= unsigned(din(19 downto  16) & "00");
            -- converted to bytes from words
          else
            hdr_length <= hdr_length;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Store the version
    --    IPv4 = 0x4
    ---------------------------------------------------------------------------
    ETHERNET_VERSION_REG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          version <= (others => '0');
        else
          if store_version = '1' then
            version <= din(23 downto  20);
          else
            version <= version;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Counter used for micsellaneous functions in the FSM
    ---------------------------------------------------------------------------
    ETHERNET_HEADER_CNT: process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_hdr_cnt = '1' then
          hdr_cnt <= (others => '0');
        else
          if en_ipv4_hdr_cnt  = '1' or en_pcol_hdr_cnt = '1' then
            hdr_cnt <= hdr_cnt + 1;
          else
            hdr_cnt <= hdr_cnt;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  For TCP length for the Pseudo header
    --    At calc_frm_length, din_big_end contains the total length of
    --      the packet starting from the IPv4 header to the end of the packet.
    --      Subtract off the IPv4 Header Length (should be 5 words / 20 bytes
    --      to get the TCP Length for the pseudo header
    ---------------------------------------------------------------------------
    ETHERNET_FRAME_LENGTH: process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          frm_length <= (others => '0');
        else
          if calc_frm_length = '1' then
          -- This is asserted for both TCP and UDP
          -- This is stored BIG Endian
            frm_length <= std_logic_vector(unsigned(din_big_end(0 to 15)) - hdr_length);
          else
            frm_length <= frm_length;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Store this information for the Pseudo Header
    --    Pseudo Header:   ________________________________
    --              Wd 0  |______ IP Source Address ______|
    --              Wd 1  |___ IP Destination Address ____|
    --              Wd 2  |__ 0 __|_PCOL _|_ TCP Length __|
    --
    ---------------------------------------------------------------------------
    ETHERNET_SA0: process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          sa0 <= (others => '0');
        else
          if store_sa_da = '1' and hdr_cnt = "011" then
            sa0 <= din(31 downto 16);
          else
            sa0 <= sa0;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Store this information for the Pseudo Header
    --    Pseudo Header:   ________________________________
    --              Wd 0  |______ IP Source Address ______|
    --              Wd 1  |___ IP Destination Address ____|
    --              Wd 2  |__ 0 __|_PCOL _|_ TCP Length __|
    --
    ---------------------------------------------------------------------------
    ETHERNET_SA1_DA0: process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          sa1 <= (others => '0');
          da0 <= (others => '0');
        else
          if store_sa_da = '1' and hdr_cnt = "100" then
            sa1 <= din(15 downto  0);
            da0 <= din(31 downto 16);
          else
            sa1 <= sa1;
            da0 <= da0;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Store this information for the Pseudo Header which is 32-bits x 3 deep
    --    Pseudo Header:   ________________________________
    --              Wd 0  |______ IP Source Address ______|
    --              Wd 1  |___ IP Destination Address ____|
    --              Wd 2  |__ 0 __|_PCOL _|_ TCP Length __|
    --
    ---------------------------------------------------------------------------
    ETHERNET_DA_HALF: process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          da1 <= (others => '0');
        else
          if store_sa_da = '1' and hdr_cnt = "000" then
            da1 <= din(15 downto  0);
          else
            da1 <= da1;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Set and hold the Pseudo Header information
    --    Big Endian Pseudo Header:    ________________________________
    --                          Wd 0  |______ IP Source Address ______|
    --                          Wd 1  |___ IP Destination Address ____|
    --                          Wd 2  |__ 0 __|_PCOL _|_ TCP Length __|
    --                  Wd 2 Example {| 0x00  | 0x06  | 0x01  | 0xFF  | }
    --
    --    Little Endian Pseudo Header: ________________________________
    --                          Wd 0  |______ IP Source Address ______|
    --                          Wd 1  |___ IP Destination Address ____|
    --                          Wd 2  |_ TCP Length __|_PCOL _|__ 0 __|
    --                  Wd 2 Example {| 0xFF  | 0x01  | 0x06  | 0x00  | }
    --
    --
    ---------------------------------------------------------------------------
    PSEUDO_HDR_WD2 : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          pseudo_data        <= (others => '0');
        else
          if tcp_ptcl_int = '1' then
          --  put back to little endian before write to BRAM
            pseudo_data       <= frm_length(8 to 15) & frm_length(0 to 7) &  X"06" & X"00";
          elsif udp_ptcl_int = '1' and calc_frm_length = '1' then
            pseudo_data       <= din(31 downto 16) & X"11" & X"00";
          else
            pseudo_data       <= pseudo_data;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  At the end of the packet, mux in the Pseudo data Wd 2 to be calculated
    --  in the CSUM.  The CSUM Actually starts with IP Source Address,
    --  but adds this word in last.
    --
    --  This is done last for commanality between TCP and UDP, since for UDP
    --  the Length is provided in the UDP Header which occurs after the CSUM
    --  starts.  In both TCP and UDP the CSUM starts at the IP Source Address
    --    Pseudo Header:   ________________________________
    --              Wd 0  |______ IP Source Address ______|
    --              Wd 1  |___ IP Destination Address ____|
    --              Wd 2  |__ 0 __|_PCOL _|_ TCP Length __|
    --
    ---------------------------------------------------------------------------
    CMB_CSUM_DIN_MUX : process (add_psdo_wd_int,pseudo_data,din,not_tcp_udp_int)
    begin

      if add_psdo_wd_int = '1' and not_tcp_udp_int = '0' then
        csum_din <= pseudo_data;
      else
        csum_din <= din;
      end if;
    end process;


    ---------------------------------------------------------------------------
    --  Set the Ethernet II flag indicator which is used to determine if
    --  the Full CSUM will be calculated.
    ---------------------------------------------------------------------------
    ETHERNET_II_REG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          eth2 <= '0';
        else
          if set_eth2 = '1' then
            eth2 <= '1';
          else
            eth2 <= eth2;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Set the Subnetwork Access Protocol (SNAP) Frame flag indicator which
    --  is used to determine if the Full CSUM will be calculated.
    ---------------------------------------------------------------------------
    ETHERNET_SNAP_REG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          snap_hit <= '0';
        else
          if set_snap = '1' then
            snap_hit <= '1';
          else
            snap_hit <= snap_hit;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Set the SNAP Frame Organizationally Unique Identifier (OUI) flag
    --  indicator which is used to determine if the Full CSUM will be
    --  calculated.
    ---------------------------------------------------------------------------
    ETHERNET_SNAP_OUI_REG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          oui_hit <= '0';
        else
          if set_oui_hit = '1' then
            oui_hit <= '1';
          else
            oui_hit <= oui_hit;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Set the VLAN flag indicator which is used to determine if the Full
    --  CSUM will be calculated.
    ---------------------------------------------------------------------------
    ETHERNET_VLAN_REG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          vlan <= '0';
        else
          if set_vlan = '1' then
            vlan <= '1';
          else
            vlan <= vlan;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Set the IPv4 protocol flag indicator which is used to determine if the
    --  Full CSUM will be calculated.
    ---------------------------------------------------------------------------
    ETHERNET_IPV4_REG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          ipv4 <= '0';
        else
          if set_ipv4 = '1' then
            ipv4 <= '1';
          else
            ipv4 <= ipv4;
          end if;
        end if;
      end if;
    end process;


    ---------------------------------------------------------------------------
    --  Set the enable to write the IPv4 header CSUM when it is time.
    ---------------------------------------------------------------------------
    DO_IPV4_HEADER : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          do_ipv4_int <= '0';
        else
          if set_ipv4hdr_only = '1' then --or do_full_csum_int = '1' then
            do_ipv4_int <= '1';
          else
            do_ipv4_int <= do_ipv4_int;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Set flag to do IPv4 header csum even though there is not a tcp or udp
    --  protocol
    ---------------------------------------------------------------------------
    IPV4_HDRCSUM_NO_PTCL : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          not_tcp_udp_int <= '0';
        elsif set_not_tcp_udp = '1' then
          not_tcp_udp_int <= '1';
        else
          not_tcp_udp_int <= not_tcp_udp_int;
        end if;
      end if;
    end process;


    ---------------------------------------------------------------------------
    --  Set the TCP protocol flag indicator which is used to determine if the
    --  Full CSUM will be calculated.
    ---------------------------------------------------------------------------
    ETHERNET_TCP_REG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          tcp_ptcl_int <= '0';
        else
          if set_ptcl = '1' and din(31 downto 24) = X"06" then
            tcp_ptcl_int <= '1';
          else
            tcp_ptcl_int <= tcp_ptcl_int;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Set the UDP protocol flag indicator which is used to determine if the
    --  Full CSUM will be calculated.
    ---------------------------------------------------------------------------
    ETHERNET_UDP_REG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          udp_ptcl_int <= '0';
        else
          if set_ptcl = '1' and din(31 downto  24) = X"11" then
            udp_ptcl_int <= '1';
          else
            udp_ptcl_int <= udp_ptcl_int;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Set the Fragment flag indicator which is used to determine if the
    --  Full CSUM will be calculated.
    --    Fragment currrently are not supported
    ---------------------------------------------------------------------------
    ETHERNET_FRAGMENT : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          fragment <= '0';
        else
          if set_fragment = '1' then
            fragment <= '1';
          else
            fragment <= fragment;
          end if;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Indicates all of the conditions were not met to perform the CSUM
    ---------------------------------------------------------------------------
--    ABORT_CHECKSUM : process(AXI_STR_TXD_ACLK)
--    begin

--      if rising_edge(AXI_STR_TXD_ACLK) then
        abort_csum <= abort_csum_int;
--      end if;
--    end process;



    ---------------------------------------------------------------------------
    --  Calculate the IPv4 Header CSUM address offsets
    --    Numerous flags are used to determine the offset
    --    Also set the BRAM write enable appropriately
    ---------------------------------------------------------------------------
    CSUM_IPV4HDR_ADDR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          csum_ipv4_hdr_addr_int <= (others => '0');
          csum_ipv4_hdr_we_int   <= (others => '0');
        elsif clr_hdr_cnt = '1' and store_sa_da = '1' and ipv4 = '1' then
          if vlan = '1' and eth2 = '1' then
            csum_ipv4_hdr_addr_int <= unsigned(csum_strt_addr) + 7;
            csum_ipv4_hdr_we_int   <= "0011";
          elsif vlan = '1' and snap_hit = '1' and oui_hit = '1' then
            csum_ipv4_hdr_addr_int <= unsigned(csum_strt_addr) + 9;
            csum_ipv4_hdr_we_int   <= "0011";
          elsif vlan = '0' and eth2 = '1' then
            csum_ipv4_hdr_addr_int <= unsigned(csum_strt_addr) + 6;
            csum_ipv4_hdr_we_int   <= "0011";
          elsif vlan = '0' and snap_hit = '1' and oui_hit = '1' then
            csum_ipv4_hdr_addr_int <= unsigned(csum_strt_addr) + 8;
            csum_ipv4_hdr_we_int   <= "0011";
          else
            csum_ipv4_hdr_addr_int <= csum_ipv4_hdr_addr_int;
            csum_ipv4_hdr_we_int   <= csum_ipv4_hdr_we_int;
          end if;
        else
          csum_ipv4_hdr_addr_int <= csum_ipv4_hdr_addr_int;
          csum_ipv4_hdr_we_int   <= csum_ipv4_hdr_we_int;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Calculate the IPv4 TCP/UDP CSUM address offsets
    --    Numerous flags are used to determine the offset
    --    Also set the BRAM write enable appropriately
    ---------------------------------------------------------------------------
    CSUM_IPV4PTCL_ADDR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_csums_int = '1' then
          do_full_csum_int       <= '0';
          csum_ptcl_addr_int     <= (others => '0');
          csum_ptcl_we_int       <= (others => '0');
        elsif clr_hdr_cnt = '1' and store_sa_da = '1' and ipv4 = '1' then
          if vlan = '1' and eth2 = '1' and tcp_ptcl_int = '1' and
             fragment = '0' then
            do_full_csum_int       <= '1';
            csum_ptcl_addr_int     <= unsigned(csum_strt_addr) + 13;
            csum_ptcl_we_int       <= "1100";
          elsif vlan = '1' and eth2 = '1' and udp_ptcl_int = '1' and
                fragment = '0' then
            do_full_csum_int       <= '1';
            csum_ptcl_addr_int     <= unsigned(csum_strt_addr) + 11;
            csum_ptcl_we_int       <= "0011";
          elsif vlan = '1' and snap_hit = '1' and oui_hit = '1' and tcp_ptcl_int = '1' and
                fragment = '0' then
            do_full_csum_int       <= '1';
            csum_ptcl_addr_int     <= unsigned(csum_strt_addr) + 15;
            csum_ptcl_we_int       <= "1100";
          elsif vlan = '1' and snap_hit = '1' and oui_hit = '1' and udp_ptcl_int = '1' and
                fragment = '0' then
            do_full_csum_int       <= '1';
            csum_ptcl_addr_int     <= unsigned(csum_strt_addr) + 13;
            csum_ptcl_we_int       <= "0011";
          elsif vlan = '0' and eth2 = '1' and tcp_ptcl_int = '1' and
                fragment = '0' then
            do_full_csum_int       <= '1';
            csum_ptcl_addr_int     <= unsigned(csum_strt_addr) + 12;
            csum_ptcl_we_int       <= "1100";
          elsif vlan = '0' and eth2 = '1' and udp_ptcl_int = '1' and
                fragment = '0' then
            do_full_csum_int       <= '1';
            csum_ptcl_addr_int     <= unsigned(csum_strt_addr) + 10;
            csum_ptcl_we_int       <= "0011";
          elsif vlan = '0' and snap_hit = '1' and oui_hit = '1' and tcp_ptcl_int = '1' and
                fragment = '0' then
            do_full_csum_int       <= '1';
            csum_ptcl_addr_int     <= unsigned(csum_strt_addr) + 14;
            csum_ptcl_we_int       <= "1100";
          elsif vlan = '0' and snap_hit = '1' and oui_hit = '1' and udp_ptcl_int = '1' and
                fragment = '0' then
            do_full_csum_int       <= '1';
            csum_ptcl_addr_int     <= unsigned(csum_strt_addr) + 12;
            csum_ptcl_we_int       <= "0011";
          else
            do_full_csum_int       <= do_full_csum_int;
            csum_ptcl_addr_int     <= csum_ptcl_addr_int;
            csum_ptcl_we_int       <= csum_ptcl_we_int;
          end if;
        else
          do_full_csum_int       <= do_full_csum_int;
          csum_ptcl_addr_int     <= csum_ptcl_addr_int;
          csum_ptcl_we_int       <= csum_ptcl_we_int;
        end if;
      end if;
    end process;


end rtl;


-------------------------------------------------------------------------------
-- tx_csum_full_calc_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_csum_full_calc_if.vhd
-- Version:         v1.00a
-- Description:     top level of embedded ip Ethernet MAC interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--                    tx_axistream_if.vhd
--                      tx_basic_if.vhd
--                      tx_csum_if.vhd
--                        tx_csum_full_if.vhd
--                          tx_csum_full_fsm.vhd
--          ->              tx_csum_full_calc_if.vhd
--                        tx_partial_csum_if.vhd
--                          tx_csum_partial_calc_if.vhd
--                      tx_vlan_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     09/16/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tx_if_pack.all;



-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------


entity tx_csum_full_calc_if is
  generic (
    -- 0 = calculate the TCP/UDP CSUM
    -- 1 = calculate the IPv4 Header CSUM
    C_IPV4_HEADER_CSUM  : integer range 0 to 1 := 0
  );
  port (
    clk               : in  std_logic;                      --  clk
    reset             : in  std_logic;                      --  reset
    clr_csums         : in  std_logic;                      --  clear the csum
    txd_tlast         : in  std_logic;                      --  axi_str_txd_tlast_dly0,
    csum_calc_en      : in  std_logic;                      --  axi_str_txd_tvalid_dly0 and axi_str_txd_tready_int_dly;

    tcp_ptcl          : in  std_logic;                      --  tcp protocol flag
    udp_ptcl          : in  std_logic;                      --  udp protocol flag
    do_ipv4hdr        : in  std_logic;                      --  only do the ipv4 header csum
    not_tcp_udp       : in  std_logic;                      --  only do the ipv4 header csum after received tlast in ptcol header
    do_full_csum      : in  std_logic;                      --  do IPv4 Ethernet II or SNAP CSUM

    do_csum           : in  std_logic;                      --  Full CSUM FLAG is set
    csum_en_b32       : in  std_logic_vector(1 downto 0);   --  enables for either IPv4 header or TCP/UDP CSUM calc bytes 3,2
    csum_en_b10       : in  std_logic_vector(1 downto 0);   --  enables for either IPv4 header or TCP/UDP CSUM calc bytes 1,0
    zeroes_en         : in  std_logic_vector(1 downto 0);   --  zeroes for either IPv4 header or TCP/UDP CSUM calc

    data_last         : in  std_logic;                      --  last data to be included in the csum calculation
    inc_txd_addr_one  : in  std_logic;                       --  increments the Tx Data Memory Address at end of a packet
    inc_txd_addr_one_early : in  std_logic;                 --  Pulses onle clock cycle early when do_csum is enabled with
                                                            --  txd_tlast and csum_calc_en

    csum_din          : in  std_logic_vector(31 downto 0);  --  Data for CSUM calculation
    csum_dout         : out std_logic_vector(15 downto 0);  --  Computed CSUM Result
    csum_we           : out std_logic_vector( 3 downto 0);  --  Tx Data Memory Write Enables to perform 16-bit write
    csum_cmplt        : out std_logic                       --  CSUM Calculation has completed
  );

end tx_csum_full_calc_if;

architecture rtl of tx_csum_full_calc_if is

  signal csum_3_2      : unsigned(16 downto 0);
  signal csum_1_0      : unsigned(16 downto 0);
  signal data_last_dly : std_logic_vector( 3 downto 0);
  signal hold          : std_logic;
  signal force_dly     : std_logic;

  begin
    -----------------------------------------------------------------------
    --  It takes additional clocks after data_last for the csum
    --  calculation to complete
    -----------------------------------------------------------------------
    CSUM_ENABLE_DELAYS : process(clk)
    begin

      if rising_edge(clk) then
        if reset = '1' or clr_csums = '1' then
          data_last_dly <= (others => '0');
        else
          data_last_dly(0)          <= data_last;
          data_last_dly(3 downto 1) <= data_last_dly(2 downto 0);
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------
    --  Calculate the 16 bit CSUM for AXI_STR_TXD_TDATA(31 downto 16)
    --    (bytes 3 and 2)
    --    This 16 bits is for the TCP csum
    -----------------------------------------------------------------------
    BYTE_3_2_CSUM : process(clk)
    begin

      if rising_edge(clk) then
        if reset = '1' or clr_csums = '1' then
          csum_3_2 <= (others => '0');
        else
          if data_last_dly(0) = '1' then
          --  add the carry at the end of the csum calculation
             csum_3_2 <= ('0' & csum_3_2(15 downto 0)) + (X"0000" & csum_3_2(16));
          elsif csum_en_b32 = "01" then
          --  continually calculate the csum for each 16 bits written to memory
            csum_3_2 <= ('0' & csum_3_2(15 downto 0)) +                  -- always zero out the carry and add the curren CSUM value to the next data
                        unsigned("000000000" & csum_din(23 downto 16)) + -- add the data to the csum
                        (X"0000" & csum_3_2(16));                        -- add the carry when it occurs


          elsif csum_en_b32 = "11" and zeroes_en(1) = '0' then
          --  when zeroes_en(1) = 1 then do not do CSUM; this is equivalent to muxing in zeroes when doing the TCP data csum calculation
          --  continually calculate the csum for each 16 bits written to memory
            csum_3_2 <= ('0' & csum_3_2(15 downto 0)) +          -- always zero out the carry and add the curren CSUM value to the next data
                        unsigned('0' & csum_din(31 downto 16)) + -- add the data to the csum
                        (X"0000" & csum_3_2(16));                -- add the carry when it occurs
          else --also handles the case when data_last = 1 and csum_en_b32 = "00" (axi_str_txd_strb = "0011" or "0001")
            csum_3_2 <= csum_3_2;
          end if;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------
    --  Calculate the 16 bit CSUM for AXI_STR_TXD_TDATA(15 downto 0)
    --    (bytes 1 and 0)
    --    This 16 bits is for either the IPv4 header csum or the UDP csum
    -----------------------------------------------------------------------
    BYTE_1_0_CSUM : process(clk)
    begin

      if rising_edge(clk) then
        if reset = '1' or clr_csums = '1' then
          csum_1_0 <= (others => '0');
        else
          if data_last_dly(1) = '1' then
          --  Both csum_3_2 and csum_1_0 are calculated, but they need to be added
          --    to each other and then checked for overflow (inc_txd_addr_one_dly2)
             csum_1_0 <= '0' & csum_3_2(15 downto 0) + csum_1_0(15 downto 0);
          elsif data_last_dly(0) = '1' or data_last_dly(2) = '1' then
          --  add the carry at the end of the data written to memory or
          --  add the carry at the end of the csum calculation
          --    (after csum 3_2 has been added to csum(1_0))
             csum_1_0 <= ('0' & csum_1_0(15 downto 0)) + (X"0000" & csum_1_0(16));
          elsif csum_en_b10 = "01" then
            --  continually calculate the csum for each 16 bits written to memory
              csum_1_0 <= ('0' & csum_1_0(15 downto 0)) +                 -- always zero out the carry and add the curren CSUM value to the next data
                          unsigned("000000000" & csum_din(7 downto  0)) + -- add the data to the csum
                          (X"0000" & csum_1_0(16));                       -- add the carry when it occurs

          elsif csum_en_b10 = "11" and zeroes_en(0) = '0' then
          --  when zeroes_en(0) = 1 then do not do CSUM; this is equivalent to muxing in zeroes when doing the ipv4 header csum calculation
          --  or when doing the UDP data csum calculation

          -- also handles when data_last = 1 (csum_en_b10 must always be 11 or 01 when null strobes are not supported)
          -- (axi_str_txd_strb = "1111" or "0111" or "0011" or "0001")
            --  when zeroes_en(0) = 1 then do not do CSUM; this is equivalent to muxing in zeroes when doing the data csum calculation
            --  continually calculate the csum for each 16 bits written to memory
            csum_1_0 <= ('0' & csum_1_0(15 downto 0)) +          -- always zero out the carry and add the curren CSUM value to the next data
                        unsigned('0' & csum_din(15 downto  0)) + -- add the data to the csum
                        (X"0000" & csum_1_0(16));                -- add the carry when it occurs
          else
            csum_1_0 <= csum_1_0;
          end if;
        end if;
      end if;
    end process;



      HOLD_REGISTER : process(clk)
      begin

        if rising_edge(clk) then
          if reset = '1' or clr_csums = '1' then
            hold     <= '0';
          else
            if (inc_txd_addr_one = '1' and (do_ipv4hdr = '1' or do_full_csum = '1') and not_tcp_udp = '0') then
            --  header CSUM or TCP/UDP CSUM is being done
              hold <= '1';
            elsif (inc_txd_addr_one = '1' and (do_ipv4hdr = '0' and do_full_csum = '0') and not_tcp_udp = '0' and do_csum = '1') then
            --  no header and no TCP/UDP CSUMs (>= 64bytes)
              hold <= '1';
            elsif (not_tcp_udp = '1' and data_last_dly(2) = '1' and inc_txd_addr_one_early = '0') or force_dly = '1' then
            --  no header and no TCP/UDP CSUMs (<64 bytes)
            --  inc_txd_addr_one cannot occure with hdr_csum_wr so use force_dly  to delay  hdr_csum_wr
              hold <= '1';
            else
              hold <= hold;
            end if;
          end if;
        end if;
      end process;


      -------------------------------------------------------------------------
      --  For packets <64 bytes when hdr_csum_wr cannot occur with inc_txd_addr_one
      -------------------------------------------------------------------------
      FORCE_DELAY : process(clk)
      begin

        if rising_edge(clk) then
          if not_tcp_udp = '1' and data_last_dly(2) = '1' and inc_txd_addr_one_early = '1' then
            force_dly <= '1';
          else
            force_dly <= '0';
          end if;
        end if;
      end process;



    -------------------------------------------------------------------------
    --  Generate the logic for the TCP/UDP CSUM
    -------------------------------------------------------------------------
    GEN_IPV4_DATA_CSUM : if C_IPV4_HEADER_CSUM = 0 generate
    begin

      --  The requirement for checksum is to invert the final value, if it is UDP and "0x0000" then
      --  set it back to "0xFFFF".  To save a step of inversion, just check it to see if it is
      --  0xFFFF before the inversion, and if it is, then do not invert it.

        csum_dout  <= x"FFFF" when (udp_ptcl = '1' and data_last_dly(3) = '1' and csum_1_0 = x"FFFF") else
                      not std_logic_vector(csum_1_0(15 downto 0));

        csum_we    <= "1100" when data_last_dly(3) = '1' and tcp_ptcl = '1' else
                      "0011" when data_last_dly(3) = '1' and udp_ptcl = '0' else
                      "0000";

        --csum_cmplt <= data_last_dly(3);





        CSUM_COMPLETE : process(clk)
        begin

          if rising_edge(clk) then
            if reset = '1' then
              csum_cmplt <= '0';
            else
              if do_csum = '1' and do_full_csum = '1' then  --did
                if data_last_dly(2) = '1' and do_full_csum = '1' then
                --  this will happen simultaneously with data_last_dly(3) when performing the csum
                  csum_cmplt <= '1';
                else
                  csum_cmplt <= '0';
                end if;
              elsif not_tcp_udp = '1' then
                if data_last_dly(0) = '1' then
                --  Not doing TCP or UDP CSUM and data ends during TCP/UDP bytes (data ends first byte after IPv4 header)
                --  delay the txd Write FSM in tx_csum_full_if until the ipv4 header is complete
                  csum_cmplt <= '1';
                else
                  csum_cmplt <= '0';
                end if;
              elsif not_tcp_udp = '0' then
                if (inc_txd_addr_one = '1' and do_ipv4hdr = '1' and do_full_csum = '0') or -- only do IPv4 header csum
                    data_last_dly(0) = '1' then -- not doing any csum, but need to set enable to exit FSMs
                  csum_cmplt <= '1';
                else
                  csum_cmplt <= '0';
                end if;
              else
                csum_cmplt <= '0';
              end if;

            end if;
          end if;
        end process;

    end generate GEN_IPV4_DATA_CSUM;

    -------------------------------------------------------------------------
    --  Generate the logic for the IPv4 Header CSUM
    -------------------------------------------------------------------------
    GEN_IPV4_HEADER_CSUM : if C_IPV4_HEADER_CSUM = 1 generate
    begin


--      HOLD_REGISTER : process(clk)
--      begin
--
--        if rising_edge(clk) then
--          if reset = '1' or clr_csums = '1' then
--            hold <= '0';
--          else
--            if inc_txd_addr_one = '1' and do_ipv4hdr = '1' then
--              hold <= '1';
--            else
--              hold <= hold;
--            end if;
--          end if;
--        end if;
--      end process;
--
      --  The requirement for checksum is to invert the final value
        csum_dout  <= not std_logic_vector(csum_1_0(15 downto 0));
        csum_we    <= "0011" when hold = '1' else
                      "0000";
        csum_cmplt <= hold;

    end generate GEN_IPV4_HEADER_CSUM;

end rtl;





-------------------------------------------------------------------------------
-- tx_csum_partial_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_csum_partial_if.vhd
-- Version:         v1.00a
-- Description:     embedded ip AXI Stream transmit interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--                    tx_axistream_if.vhd
--                      tx_basic_if.vhd
--                      tx_csum_if.vhd
--                        tx_csum_full_if.vhd
--                          tx_csum_full_fsm.vhd
--                          tx_csum_full_calc_if.vhd
--          ->            tx_csum_partial_if.vhd
--                          tx_csum_partial_calc_if.vhd
--                      tx_vlan_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tx_if_pack.all;

-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity tx_csum_partial_if is
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data


    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0)   --  Tx AXI-Stream Control to Memory Full Flag

  );

end tx_csum_partial_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of tx_csum_partial_if is


-------------------------------------------------------------------------------
--  Start Partial CSUM
-------------------------------------------------------------------------------
  constant zeroes_txc                     : std_logic_vector(c_TxC_write_width_b -1 downto c_TxC_addrb_width) := (others => '0');
  constant zeroes_txd                     : std_logic_vector(c_TxC_write_width_b -1 downto c_TxD_addrb_width) := (others => '0');
  constant zeroes_txd_2                   : std_logic_vector(c_TxC_write_width_b -1 downto c_TxD_addrb_width + 2 ) := (others => '0');

  type TXC_WR_FSM_TYPE is (
                       TXC_ADDR2_WR,
                       TXC_ADDR0_WR,
                       WAIT_WR_CMPLT,
                       TXC_WD0,
--                       WAIT_TXD_FULL,
                       TXC_WD1,
                       WAIT_ADDR2_COMPARE_CMPLT,--added for BRAM async clocks
                       TXC_WD2,
                       TXC_WD3,
                       TXC_WD4,
                       WAIT_ADDR0_COMPARE_CMPLT,--added for BRAM async clocks
                       TXC_WD5,
                       WAIT_TXD_CMPLT,
                       WAIT_TXD_MEM,
                       WR_TXC_PNTR,
                       WAIT_CSUM_END,
                       WR_TXD_END_PNTR
                      );
  signal txc_wr_cs, txc_wr_ns             : TXC_WR_FSM_TYPE;

  type TXD_WR_FSM_TYPE is (
                       IDLE,
                       TXD_PRM,
                       TXD_WRT,
                       MEM_FULL,
                       CLR_FULL,
                       WAIT_WR1,
                       WAIT_WR2,
                       WAIT_CSUM,
                       WAIT_COMPARE_CMPLT
                      );
  signal txd_wr_cs, txd_wr_ns             : TXD_WR_FSM_TYPE;

  signal txc_min_wr_addr                  : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_rsvd_wr_addr                 : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_max_wr_addr                  : std_logic_vector(c_TxC_addrb_width -1 downto 0);

  signal txc_wr_addr0                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr1                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr2                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr3                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr5                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr6                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);

  signal axi_str_txc_tready_int           : std_logic;
  signal axi_str_txc_tready_int_dly       : std_logic;
  signal axi_str_txc_tvalid_dly0          : std_logic;
  signal axi_str_txc_tlast_dly0           : std_logic;
--  signal axi_str_txc_tstrb_dly0           : std_logic_vector(3 downto 0);
  signal axi_str_txc_tdata_dly0           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal clr_txc_trdy                     : std_logic;

  signal axi_str_txd_tready_int           : std_logic;
  signal axi_str_txd_tready_int_dly       : std_logic;
  signal axi_str_txd_tvalid_dly0          : std_logic;
  signal axi_str_txd_tlast_dly0           : std_logic;
  signal axi_str_txd_tstrb_dly0           : std_logic_vector(3 downto 0);
  signal axi_str_txd_tdata_dly0           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal axi_str_txd_tdata_dly1           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal clr_txd_trdy                     : std_logic;

  signal set_txc_addr_0                   : std_logic;
  signal txc_addr_0_dly1                  : std_logic;
  signal txc_addr_0_dly2                  : std_logic;
  signal set_txc_addr_1                   : std_logic;
  signal txc_addr_1                       : std_logic;
  signal set_txc_addr_2                   : std_logic;
  signal txc_addr_2                       : std_logic;
  signal set_txc_addr_4_n                 : std_logic;
  signal set_txc_addr_3                   : std_logic;
  signal clr_txc_addr_3                   : std_logic;
  signal txc_addr_3_dly                   : std_logic;
  signal txc_addr_3_dly2                  : std_logic;
  signal txc_addr_3_dly3                  : std_logic;
  signal inc_txd_addr_one                 : std_logic;
  signal set_txc_trdy                     : std_logic;
  signal set_txc_trdy2                    : std_logic;
  signal clr_txc_trdy2                    : std_logic;
  signal set_txcwr_rd_addr                : std_logic;
  signal set_txcwr_wr_end                 : std_logic;
  signal set_txc_en                       : std_logic;
  signal set_txc_we                       : std_logic;
  signal txc_we                           : std_logic;
  signal txc_we_dly1                      : std_logic;
  signal txc_we_dly2                      : std_logic;

  signal addr_2_en                        : std_logic;
  signal addr_2_en_dly1                   : std_logic;
  signal addr_2_en_dly2                   : std_logic;

  signal txc_mem_full                     : std_logic;
  signal txc_mem_not_full                 : std_logic;
  signal txc_mem_afull                    : std_logic;
  signal txc_mem_wr_addr                  : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_0                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_1                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_last             : std_logic_vector(c_TxC_addrb_width   -1 downto 0);

  signal Axi_Str_TxC_2_Mem_Addr_int       : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal Axi_Str_TxC_2_Mem_We_int         : std_logic_vector(0 downto 0);
  signal txc_mem_wr_addr_plus1            : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_plus2            : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_rd_addr2_pntr                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_rd_addr2_pntr_1              : std_logic_vector(c_TxC_addrb_width   -1 downto 0);


  -- Set to the full width of the write data bus
  signal Axi_Str_TxC_2_Mem_Din_int        : std_logic_vector(c_TxC_write_width_b -1 downto 0);

  signal set_axi_flag                     : std_logic;
  signal set_csum_cntrl                   : std_logic;
  signal set_csum_begin_insert            : std_logic;
  signal set_csum_rsvd_init               : std_logic;
  signal axi_flag                         : std_logic_vector( 3 downto 0);
  signal csum_cntrl                       : std_logic_vector( 1 downto 0);

  signal set_first_packet                 : std_logic;
  signal wrote_first_packet               : std_logic;
  signal inc_txd_wr_addr                  : std_logic;
  signal set_txd_we                       : std_logic_vector( 3 downto 0);
  signal set_txd_en                       : std_logic;
  signal set_txd_rdy                      : std_logic;
  signal clr_txd_rdy                      : std_logic;
  signal clr_full_pntr                    : std_logic;
  signal halt_pntr_update                 : std_logic;
  signal disable_txd_trdy                 : std_logic;
  signal disable_txd_trdy_dly             : std_logic;
  signal disable_txc_trdy                 : std_logic;
  signal disable_txc_trdy_dly             : std_logic;

  signal txd_rdy                          : std_logic;
  signal axi_str_txd_2_mem_addr_int       : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_last  : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_mins1 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus1 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus2 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus3 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus4 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txd_mem_full                     : std_logic;
  signal txd_mem_not_full                 : std_logic;
  signal txd_mem_afull                    : std_logic;
  signal axi_str_txd_2_mem_we_int         : std_logic_vector( 3 downto 0);
  signal axi_str_txd_2_mem_en_int         : std_logic;

  signal txd_rd_pntr                      : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_1                    : std_logic_vector(c_TxD_addrb_width -1 downto 0);

  signal txd_min_wr_addr                  : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_max_wr_addr                  : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_max_wr_addr_minus4           : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_hold_plus3           : std_logic_vector(c_TxD_addrb_width -1 downto 0);

  signal txd_rd_pntr_hold                 : std_logic_vector(c_TxD_addrb_width -1 downto 0);

  signal csum_begin_int                   : std_logic_vector(15 downto 0);
  signal csum_begin                       : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal csum_begin_bytes                 : std_logic_vector( 1 downto 0);
  signal csum_insert_int                  : std_logic_vector(15 downto 0);
  signal csum_insert                      : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal csum_insert_bytes                : std_logic_vector( 1 downto 0);
  signal csum_init                        : std_logic_vector(15 downto 0);

  constant zeroes_csum                    : std_logic_vector(15 downto c_TxD_addrb_width) := (others => '0');

  signal load_csum_int                    : std_logic;
  signal csum_addr                        : std_logic_vector(c_TxD_addrb_width   -1 downto 0);


  signal do_csum                          : std_logic;
  signal csum_result                      : std_logic_vector(15 downto 0);
  signal csum_en                          : std_logic;
  signal csum_we                          : std_logic_vector(3 downto 0);

  signal csum_en_dly                      : std_logic;
  signal csum_cmplt                       : std_logic;

  signal tx_init_in_prog_int              : std_logic;
  signal init_bram                        : std_logic;

  signal txc_rd_addr0                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txc_rd_addr2                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txc_rd_addr3                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);

  signal set_txd_mem_full                 : std_logic;
  signal clr_txd_mem_full                 : std_logic;
  signal set_txd_mem_afull                : std_logic;

  signal compare_addr0                    : std_logic;
  signal compare_addr0_cmplt              : std_logic;

  signal compare_addr2                    : std_logic;
  signal compare_addr2_cmplt              : std_logic;
  signal compare_addr2_cmplt_dly          : std_logic;

  signal update_bram_cnt                  : unsigned(7 downto 0);

  signal enable_compare_addr0_cmplt       : std_logic;
  signal end_addr_byte_offset             : std_logic_vector(1 downto 0);


  signal check_full                       : std_logic;
  signal update_rd_pntrs                  : std_logic;


  begin

    -----------------------------------------------------------------------------
    --  The TxC BRAM is set up to to always store the current TxD Read and Write
    --    pointers in the first two locations (0x0 and 0x1) of the Memory
    --    respectivively.  The current TxC Read and write pointer are always
    --    stored in the the next two locations (0x2 and 0x3) of the Memory
    --    respectively.  The End addresses for each packet are then stored
    --    in the remaing Memory locations starting at address 0x4.  After
    --    the end pointer to the maximum address has been written, if the
    --    memory is not full, the address pointer will loop back to address
    --    0x4 and write the end pointer for the next packet.
    --
    --                                   BRAM
    --                             Write       Read
    --                           _____________________
    --                          |__________|_________| <-- TxD Rd Pointer
    --      TxD Wr Pointer -->  |__________|_________|
    --                          |__________|_________| <-- TxC Rd Pointer
    --      TxC Wr Pointer -->  |__________|_________|
    --      Packet 0 End   -->  |__________|_________|  --> Packet 0 End
    --      Packet 1 End   -->  |__________|_________|  --> Packet 1 End
    --      Packet 2 End   -->  |__________|_________|  --> Packet 2 End
    --         .                |__________|_________|         .
    --         .                |__________|_________|         .
    --         .                |__________|_________|         .
    --      Packet n End   -->  |__________|_________|  --> Packet n End
    --
    -----------------------------------------------------------------------------

    -----------------------------------------------------------------------------
    --  Create the full and empty comparison values for the S6 and V6 since
    --  1 S6 BRAM = 1/2 V6 BRAM
    -----------------------------------------------------------------------------
    GEN_TXC_MIN_MAX_WR_FLAG : for i in (c_TxC_addrb_width-1) downto 0 generate
      txc_min_wr_addr(i)  <= '1' when (i = 2)          else '0'; -- do not loop back to 0x0; loop to 0x4
      txc_max_wr_addr(i)  <= '0' when (i = 0 or i = 1) else '1';
      txc_wr_addr0(i)     <= '0';
      txc_wr_addr1(i)     <= '1' when (i = 0)          else '0';
      txc_wr_addr2(i)     <= '1' when (i = 1)          else '0';
      txc_wr_addr3(i)     <= '1' when (i = 0 or i = 1) else '0';
      txc_wr_addr5(i)     <= '1' when (i = 0 or i = 2) else '0';
      txc_wr_addr6(i)     <= '1' when (i = 1 or i = 2) else '0';
    end generate GEN_TXC_MIN_MAX_WR_FLAG;

    GEN_TXD_MIN_MAX_WR_FLAG : for i in (c_TxD_addrb_width-1) downto 0 generate
      txd_min_wr_addr(i)        <= '1' when (i = 0) else '0';
      txd_max_wr_addr_minus4(i) <= '0' when (i = 2) else '1';
      txd_max_wr_addr(i)        <= '1';
    end generate GEN_TXD_MIN_MAX_WR_FLAG;


    GEN_TXC_MIN_MAX_RD_FLAG : for i in (c_TxD_addrb_width-1) downto 0 generate
      txc_rd_addr0(i)     <= '0';
      txc_rd_addr2(i)     <= '1' when (i = 1)          else '0';
      txc_rd_addr3(i)     <= '1' when (i = 0 or i = 1) else '0';
    end generate GEN_TXC_MIN_MAX_RD_FLAG;




    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Control Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXC_CONTROL : process(AXI_STR_TXC_ACLK)
    begin
      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          axi_str_txc_tvalid_dly0 <= '0';
          axi_str_txc_tlast_dly0  <= '0';
          clr_txc_trdy           <= '0';
        else
          axi_str_txc_tvalid_dly0 <= axi_str_txc_tvalid;
          axi_str_txc_tlast_dly0  <= axi_str_txc_tlast;
          if axi_str_txc_tvalid = '1' and axi_str_txc_tlast = '1' and axi_str_txc_tready_int = '1' then
            clr_txc_trdy <= '1';
          else
            clr_txc_trdy <= '0';
          end if;
        end if;
      end if;
    end process;

    -- Register the incoming AXI Stream Control Data Bus
    -----------------------------------------------------------------------------
    REG_TXC_IN : process(AXI_STR_TXC_ACLK)
    begin
      if rising_edge(AXI_STR_TXC_ACLK) then
--          axi_str_txc_tstrb_dly0  <= axi_str_txc_tstrb;
          axi_str_txc_tdata_dly0  <= axi_str_txc_tdata;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  AXI Stream TX Control State Machine - combinational/combinatorial
    --    Used to register the incoming control and checksum information
    --    This state machine will throttle the Transmit AXI Stream Data state
    --      machine until after the control information has been received.
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXC_CMB : process (txc_wr_cs,axi_str_txc_tvalid_dly0,
      axi_str_txc_tlast_dly0,axi_str_txd_tlast_dly0,
      axi_str_txd_tvalid_dly0,txc_addr_3_dly,
      wrote_first_packet,axi_str_txc_tready_int_dly,axi_str_txd_tready_int_dly,
      disable_txd_trdy_dly,disable_txc_trdy_dly,do_csum,csum_cmplt,
      compare_addr2_cmplt,compare_addr2_cmplt_dly,compare_addr0_cmplt,
      update_bram_cnt,txc_mem_full)

    begin


      set_axi_flag           <= '0';
      set_csum_cntrl         <= '0';
      set_csum_begin_insert  <= '0';
      set_csum_rsvd_init     <= '0';
      set_txc_addr_0         <= '0';
      set_txc_addr_1         <= '0';
      set_txc_addr_2         <= '0';
      set_txc_addr_3         <= '0';
      set_txc_addr_4_n       <= '0';
      clr_txc_addr_3         <= '0';
      set_txcwr_rd_addr      <= '0';  --  sets the write side, read address to 0x0
      set_txcwr_wr_end       <= '0';  --  writes the end address to the memory in the next available location
      set_txc_en             <= '0';  --  the enable bit to the write side of the memory
      set_txc_we             <= '0';  --  the write enable bit to the write side of the memory
      inc_txd_addr_one       <= '0';
      set_txc_trdy           <= '0';
      init_bram              <= '0';
      compare_addr2          <= '0';
      compare_addr0          <= '0';
      set_txc_trdy2          <= '0';
      clr_txc_trdy2          <= '0';
      enable_compare_addr0_cmplt <= '0';

      case txc_wr_cs is
        when TXC_ADDR2_WR =>
          set_txc_addr_2         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          txc_wr_ns              <= TXC_ADDR0_WR;
        when TXC_ADDR0_WR =>
          set_txc_addr_0         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          txc_wr_ns              <= WAIT_WR_CMPLT;
        when WAIT_WR_CMPLT =>
          set_txc_addr_0         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          set_txc_trdy2          <= '1';
          txc_wr_ns              <= TXC_WD0;
        when TXC_WD0 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' and
             (wrote_first_packet = '0' or txc_addr_3_dly = '1') then
            set_txc_addr_2         <= '1';  --Set the address to get the TxC Rd Address Pointer
            set_txc_en             <= '1';
            set_axi_flag           <= '1';
            clr_txc_addr_3         <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD1;
          else
            set_txc_addr_2         <= '0';  --Set the address to get the TxC Rd Address Pointer
            set_txc_en             <= '0';
            set_axi_flag           <= '0';
            clr_txc_addr_3         <= '0';
            compare_addr2          <= '0';
            txc_wr_ns              <= TXC_WD0;
          end if;

        when TXC_WD1 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_txc_trdy2          <= '0';
            set_csum_cntrl         <= '1';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD2;--WAIT_ADDR2_COMPARE_CMPLT;
          elsif axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '0' then
          -- need to force txc trdy HIGH since TVALID throttled
            set_txc_trdy2          <= '1';
            set_csum_cntrl         <= '0';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= WAIT_ADDR2_COMPARE_CMPLT;
          else
            set_txc_trdy2          <= '0';
            set_csum_cntrl         <= '0';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD1;
          end if;

        when WAIT_ADDR2_COMPARE_CMPLT =>
        -- now clear txc trdy to only allow a one clock pulse HIGH
          clr_txc_trdy2          <= '1';
          set_txc_addr_2         <= '1';
          set_txc_en             <= '1';
          compare_addr2          <= '1';
          txc_wr_ns              <= TXC_WD1;

        when TXC_WD2 =>
        -- Txc Tready has already been disabled
        --  wait for compare_addr2_cmplt, then
        --  set_txc_trdy2 will force axi_str_txc_tready_int_dly HIGH
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_csum_begin_insert      <= '1';
            set_txc_addr_2         <= '0';
            set_txc_en             <= '0';
            compare_addr2          <= '0';
            set_txc_trdy2          <= '0';
            txc_wr_ns                  <= TXC_WD3;
          else
            if axi_str_txc_tvalid_dly0 = '0'  or
               (txc_mem_full = '1' and axi_str_txc_tvalid_dly0 = '1') then
            --  If full wait for FULL and TVALID
            --  This will allow next elsif to be hit properly
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '1';
              set_txc_en             <= '1';
              compare_addr2          <= '1';
              set_txc_trdy2          <= '0';
              txc_wr_ns              <= TXC_WD2;


            elsif axi_str_txc_tvalid_dly0 = '1' and
              (compare_addr2_cmplt = '1' or compare_addr2_cmplt_dly = '1') then
              --  when full is '0', only need compare_addr2_cmplt to set set_txc_trdy2
              --    which will then allow this state to be exited to TXD_WD3
              --  when full is '1', then will need compare_addr2_cmplt_dly to to set set_txc_trdy2
              --    which will then allow this state to be exited to TXD_WD3
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '0';
              set_txc_en             <= '0';
              compare_addr2          <= '0';
              set_txc_trdy2          <= '1';
              txc_wr_ns                  <= TXC_WD2;
            else
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '1';
              set_txc_en             <= '1';
              compare_addr2          <= '1';
              set_txc_trdy2          <= '0';
              txc_wr_ns                  <= TXC_WD2;
            end if;
          end if;
        when TXC_WD3 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
          --  This is the earliest state to check for TxC FULL from TXC_WD0 state addr_2
          --  Register data, then assert full = 2 clks from rd
          --    Not FULL so write TxC Write Pointer to addr 0x3
            set_csum_rsvd_init         <= '1';
            txc_wr_ns                  <= TXC_WD4;
          else
            set_csum_rsvd_init         <= '0';
            txc_wr_ns                  <= TXC_WD3;
          end if;
        when TXC_WD4 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_txc_addr_0             <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            txc_wr_ns                  <= TXC_WD5;
          else
            set_txc_addr_0             <= '0';  --Set the address to get the TxD Rd Address Pointer
            set_txc_en                 <= '0';
            compare_addr0              <= '0';
            txc_wr_ns                  <= TXC_WD4;
          end if;
        when TXC_WD5 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' and axi_str_txc_tlast_dly0 = '1' then
            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '1';
            txc_wr_ns                  <= WAIT_ADDR0_COMPARE_CMPLT;
          else
            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '0';
            txc_wr_ns                  <= TXC_WD5;
          end if;
        when WAIT_ADDR0_COMPARE_CMPLT =>
          if compare_addr0_cmplt = '1' then
            set_txc_addr_1             <= '1'; -- this is one clock early, so do not set the we enable yet
            set_txc_en                 <= '1';
            set_txc_we                 <= '1';

            set_txc_addr_0             <= '0';
            set_txc_en                 <= '0';
            compare_addr0              <= '0';
            enable_compare_addr0_cmplt <= '0';
            txc_wr_ns                  <= WAIT_TXD_CMPLT;
          else
            set_txc_addr_1             <= '0';
            set_txc_en                 <= '0';
            set_txc_we                 <= '0';

            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '1';
            txc_wr_ns                  <= WAIT_ADDR0_COMPARE_CMPLT;
          end if;



        when WAIT_TXD_CMPLT =>
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1'  and
             axi_str_txd_tlast_dly0 = '1' then
            set_txc_addr_0        <= '0';
            set_txc_addr_1        <= '1';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WR_TXD_END_PNTR;
          elsif disable_txd_trdy_dly = '1' then
          -- Txd mem is full so get the current read pointer
          --  This can occure after tlast so check it in the following states
            set_txc_addr_0        <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_addr_1        <= '0';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_MEM;
          elsif update_bram_cnt(7) = '1'  then
          --Writing the current TxC write pointer so the read side can monitor it
            set_txc_addr_1        <= '1';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          else
            set_txc_addr_1        <= '0'; --Writing the current TxC write pointer so the read side can monitor it
            set_txc_addr_2        <= '0';
            set_txc_en            <= '0';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          end if;
        when WAIT_TXD_MEM =>
          if disable_txd_trdy_dly = '1' then
            -- Txd mem is full so get the current read pointer
            set_txc_addr_0        <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_addr_1        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_MEM;
          else
            set_txc_addr_0        <= '0';
            set_txc_addr_1        <= '1'; -- this is one clock early, so do not set the we enable yet
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          end if;
        when WR_TXD_END_PNTR =>
          if do_csum = '1' then
            inc_txd_addr_one      <= '1';
            set_txc_addr_4_n      <= '0'; -- Write the TxC End Value to address 0x4 - 0xn
            set_txc_en            <= '0';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_CSUM_END;
          else
            inc_txd_addr_one      <= '1';
            set_txc_addr_4_n      <= '1'; -- Write the TxC End Value to address 0x4 - 0xn
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WR_TXC_PNTR;
          end if;

        when WAIT_CSUM_END =>
          if csum_cmplt = '1' then
            inc_txd_addr_one      <= '0'; -- already incremented in WR_TXC_PNTR state
            set_txc_addr_4_n      <= '1'; -- Write the TxC end pointer value to start the tx clint FSM
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WR_TXC_PNTR;
          else
            inc_txd_addr_one      <= '0'; -- already incremented in WR_TXC_PNTR state
            set_txc_addr_4_n      <= '0';
            set_txc_en            <= '0';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_CSUM_END;
          end if;

        when WR_TXC_PNTR =>
          if disable_txc_trdy_dly = '1' then
            set_txc_addr_0        <= '1';
            set_txc_addr_3        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            set_txc_trdy          <= '0';
            txc_wr_ns             <= WR_TXC_PNTR;
          else
            set_txc_addr_0        <= '0'; -- Write the TxC end pointer value to start the tx clint FSM
            set_txc_addr_3        <= '1';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            set_txc_trdy          <= '1';
            txc_wr_ns             <= TXC_WD0;
          end if;

--        when WR_TXC_PNTR =>
--            set_txc_addr_3        <= '1'; -- Write the TxC end pointer value to start the tx clint FSM
--            set_txc_addr_0        <= '0';
--            set_txc_en            <= '1';
--            set_txc_we            <= '1';
--            txc_wr_ns             <= TXC_WD0;

        when others =>
          txc_wr_ns                <= TXC_ADDR2_WR;
      end case;
    end process;

    -----------------------------------------------------------------------------
    -- AXI Stream TX Control State Machine Sequencer
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXC_SEQ : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_wr_cs <= TXC_ADDR2_WR;
        else
          txc_wr_cs <= txc_wr_ns;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    -- Delay the last write to TxC memory of the first packet after reset
    -----------------------------------------------------------------------------
    TX_INIT_INDICATOR_DLYS : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_addr_3_dly2 <= '0';
          txc_addr_3_dly3 <= '0';
        else
          txc_addr_3_dly2 <= txc_addr_3_dly;
          txc_addr_3_dly3 <= txc_addr_3_dly2;
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    -- Use above delay to hold off Tx Client FSM from starting until all
    --    TxD and TxC pointer information has been written to memory
    --
    --    This signal goes through a clock crossing circuit before it is
    --      registered in the Tx Client clock domain and used to start the
    --      Tx Client Read FSM
    -----------------------------------------------------------------------------
    TX_INIT_INDICATOR : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          tx_init_in_prog_int <= '1';
        else
          if txc_addr_3_dly3 = '1' then
            tx_init_in_prog_int <= '0';
          else
            tx_init_in_prog_int <= tx_init_in_prog_int;
          end if;
        end if;
      end if;
    end process;

    tx_init_in_prog <= tx_init_in_prog_int;

    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_1_TXD_WR_PNTR : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_1 = '1' then
          txc_addr_1 <= '1';
        else
          txc_addr_1 <= '0';
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_3_DELAY : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' or clr_txc_addr_3 = '1' then
          txc_addr_3_dly  <= '0';
        elsif set_txc_addr_3 = '1' then
          txc_addr_3_dly <= '1';
        else
          txc_addr_3_dly <= txc_addr_3_dly;
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    --  Generate address that will hold the End Address
    -----------------------------------------------------------------------------
    TXC_WR_ADDR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_mem_wr_addr      <= txc_min_wr_addr;
          txc_mem_wr_addr_last <= txc_wr_addr3;
          txc_mem_wr_addr_0    <= txc_wr_addr5;
          txc_mem_wr_addr_1    <= txc_wr_addr6;
        else
          if set_txc_addr_3 = '1' then
            --  increment the address for the next packet
            --  use the delayed signal to increment after the current address
            --  can be written
            if txc_mem_wr_addr = txc_max_wr_addr then
              --  if the max address is reached, loop to address 0x4
              txc_mem_wr_addr      <= txc_mem_wr_addr_0;
              txc_mem_wr_addr_last <= txc_wr_addr3;
              txc_mem_wr_addr_0    <= txc_mem_wr_addr_1;  --plus1
              txc_mem_wr_addr_1    <= txc_wr_addr6;       --plus2
            else
              --  otherwise just increment it
              txc_mem_wr_addr      <= txc_mem_wr_addr_0;
              txc_mem_wr_addr_last <= txc_mem_wr_addr;
              txc_mem_wr_addr_0    <= txc_mem_wr_addr_1;
              txc_mem_wr_addr_1    <= std_logic_vector(unsigned(txc_mem_wr_addr_1) + 1);
            end if;
          else -- Hold the current address until something changes
            txc_mem_wr_addr      <= txc_mem_wr_addr;
            txc_mem_wr_addr_last <= txc_mem_wr_addr_last;
            txc_mem_wr_addr_0    <= txc_mem_wr_addr_0;
            txc_mem_wr_addr_1    <= txc_mem_wr_addr_1;
          end if;
        end if;
      end if;
    end process;




    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_0_DELAY : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        txc_addr_0_dly1 <= set_txc_addr_0;
        txc_addr_0_dly2 <= txc_addr_0_dly1;
      end if;

    end process;


    -----------------------------------------------------------------------------
    --  Generate address that will hold the End Address
    -----------------------------------------------------------------------------
    MEM_TXC_WR_ADDR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then

        if set_txc_addr_4_n = '1' and set_txc_we = '1' then
          -- Provide the address for the End of packet address
          Axi_Str_TxC_2_Mem_Addr_int <= txc_mem_wr_addr;
        elsif set_txc_addr_3 = '1' and set_txc_we = '1' then
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr3; --set txc wr pointer
        elsif txc_addr_2 = '1' and  (txc_we = '0' or init_bram = '1') then
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr2; --get txc rd pointer
        elsif set_txc_addr_0 = '1' and (set_txc_we = '0' or init_bram = '1') then
          --  Monitor the read pointer for a full
          --  condition in the TxD Memory
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr0;
        elsif set_txc_addr_1 = '1' then
          --  Set the TxD write pointer to
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr1;
        else
          Axi_Str_TxC_2_Mem_Addr_int <= (others => '0');
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_Addr <= Axi_Str_TxC_2_Mem_Addr_int;
    txc_mem_wr_addr_plus1  <= txc_mem_wr_addr_0;
    txc_mem_wr_addr_plus2  <= txc_mem_wr_addr_1;

    -----------------------------------------------------------------------------
    --  This process remaps the strobe signal to the byte address offset minus
    --  one byte.
    -----------------------------------------------------------------------------
    END_ADDRESS_BYTE_OFFSET : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txD = '1' then
          end_addr_byte_offset <= (others => '0');
        elsif axi_str_txd_tlast_dly0 = '1' and axi_str_txd_tvalid_dly0 = '1' and
              axi_str_txd_tready_int_dly = '1' then
          case axi_str_txd_tstrb_dly0 is
            when "1111" => end_addr_byte_offset <= "11";
            when "0111" => end_addr_byte_offset <= "10";
            when "0011" => end_addr_byte_offset <= "01";
            when others => end_addr_byte_offset <= "00";
          end case;
        else
          end_addr_byte_offset <= end_addr_byte_offset;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_WR_ADDR_VALUE : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' or init_bram = '1' then
          Axi_Str_TxC_2_Mem_Din_int <= (others => '0');

        elsif set_txc_addr_4_n = '1' and do_csum = '0' then
        --write the ending address of the packet to memory minus one byte
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd_2 & axi_str_txd_2_mem_addr_int & end_addr_byte_offset;
        elsif set_txc_addr_4_n = '1' and do_csum = '1' then
        -- Increment already happened so use current value
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd_2 & axi_str_txd_2_mem_addr_int_mins1 & end_addr_byte_offset;
        elsif set_txc_addr_3 = '1' then
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txc & txc_mem_wr_addr;
        else
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd & axi_str_txd_2_mem_addr_int_plus1;
        end if;
      end if;
    end process;



    Axi_Str_TxC_2_Mem_Din <= Axi_Str_TxC_2_Mem_Din_int;

  --  Axi_Str_TxC_2_Mem_En  <= '1';
    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if (set_txc_en = '1' and set_txc_addr_2 = '0') or
           addr_2_en = '1' or init_bram = '1' then
          Axi_Str_TxC_2_Mem_En <= '1';
        else
          Axi_Str_TxC_2_Mem_En <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_WR_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_we = '1' then
          Axi_Str_TxC_2_Mem_We_int(0) <= '1';
        else
          Axi_Str_TxC_2_Mem_We_int(0) <= '0';
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_We <= Axi_Str_TxC_2_Mem_We_int;


    -----------------------------------------------------------------------------
    --  Delay set_txc_addr_2 to align with data
    -----------------------------------------------------------------------------
    TXC_ADDR2_DLY : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_2 = '1' then
          txc_addr_2  <= set_txc_addr_2;
        else
          txc_addr_2  <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay set_txc_we to align with address
    -----------------------------------------------------------------------------
    TXC_WE_DLY : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_we = '1' then
          txc_we  <= set_txc_we;
        else
          txc_we  <= '0';
        end if;
        txc_we_dly1 <= txc_we;
        txc_we_dly2 <= txc_we_dly1;

      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay set_txc_we to align with address
    -----------------------------------------------------------------------------
    ADDR2_MEM_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_2 = '1' and  set_txc_en = '1' then
          addr_2_en  <= set_txc_en;
        else
          addr_2_en  <= '0';
        end if;
        addr_2_en_dly1 <= addr_2_en;
        addr_2_en_dly2 <= addr_2_en_dly1;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Get the read pointer to check for FULL
    --  With ASYNC BRAM clock cannot read/write same address in memory at same
    --  time unless timing is met, so read until data matches
    -----------------------------------------------------------------------------
    MEM_TXC_RD_ADDR_PNTR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_rd_addr2_pntr_1 <= (others => '0');
          txc_rd_addr2_pntr   <= txc_min_wr_addr;
          compare_addr2_cmplt <= '0';
          compare_addr2_cmplt_dly <= '0';
        else

          if set_txc_addr_2 = '1' and addr_2_en_dly2 = '1' and txc_we_dly2 = '0' then
            txc_rd_addr2_pntr_1 <= Axi_Str_TxC_2_Mem_Dout(c_TxC_addrb_width -1 downto 0);

            if Axi_Str_TxC_2_Mem_Dout(c_TxC_addrb_width -1 downto 0) = txc_rd_addr2_pntr_1  and
               compare_addr2_cmplt = '0' then
              txc_rd_addr2_pntr   <= txc_rd_addr2_pntr_1;
              compare_addr2_cmplt <= '1';
            else
              txc_rd_addr2_pntr   <= txc_rd_addr2_pntr;
              compare_addr2_cmplt <= '0';
            end if;

          else
            txc_rd_addr2_pntr_1 <= txc_rd_addr2_pntr_1;
            txc_rd_addr2_pntr   <= txc_rd_addr2_pntr;
            compare_addr2_cmplt <= '0';
          end if;
          compare_addr2_cmplt_dly <= compare_addr2_cmplt;

        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Full flag indicator
    --    Does not begin comparison until 1st packet is written to memory
    -----------------------------------------------------------------------------
    TXC_FULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txc = '1' then
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
        elsif txc_mem_full = '1' and
           compare_addr2_cmplt = '1' and compare_addr2_cmplt_dly = '0' then
           --increments after it goes full, so use txc_mem_wr_addr for compare
          if txc_mem_wr_addr /= txc_rd_addr2_pntr then
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
          else
            txc_mem_full     <= txc_mem_full;
            txc_mem_not_full <= txc_mem_not_full;
          end if;
        elsif set_txc_addr_3 = '1' and set_txc_we = '1' then
          if txc_mem_wr_addr_plus1 = txc_rd_addr2_pntr then
            txc_mem_full     <= '1';
            txc_mem_not_full <= '0';
          else
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
          end if;
        else
          txc_mem_full     <= txc_mem_full;
          txc_mem_not_full <= txc_mem_not_full;
        end if;
      end if;
    end process;

    TXC_AFULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if txc_mem_wr_addr_plus2 = txc_rd_addr2_pntr then
          txc_mem_afull     <= '1';
        else
          txc_mem_afull     <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Throttle AXI Stream TxC
    --    Do not assert unless TxD is not in progress and the memory can
    --    accept data
    -----------------------------------------------------------------------------
    TXC_READY : process(AXI_STR_TXD_ACLK)
    begin



      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txc = '1' or clr_txc_trdy = '1' or clr_txc_trdy2 = '1' or
             set_txd_rdy = '1' or (txd_rdy = '1' and clr_txd_rdy = '0') or disable_txc_trdy = '1' or
             (AXI_STR_TXC_TLAST = '1' and AXI_STR_TXC_TVALID = '1' and axi_str_txc_tready_int = '1') or
             (compare_addr2 = '1' and axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1') then --do not need compare_addr0 because will clr at TLAST
          axi_str_txc_tready_int <= '0';
        else

          if txc_addr_3_dly = '1' then
            if (txc_mem_wr_addr = txc_rd_addr2_pntr and txc_mem_full = '1') then
              axi_str_txc_tready_int <= '0';
            elsif txc_mem_wr_addr = txc_rd_addr2_pntr and
                Axi_Str_TxC_2_Mem_We_int(0) = '1' then
              axi_str_txc_tready_int <= '0';
            else
              axi_str_txc_tready_int <= axi_str_txc_tready_int;
            end if;
          elsif set_txc_trdy = '1' then
            axi_str_txc_tready_int <= '1';
          elsif set_txc_trdy2 = '1' then
          --  need to force it high after address compare and after reset
            axi_str_txc_tready_int <= '1';
          else
            axi_str_txc_tready_int <= axi_str_txc_tready_int;
          end if;
        end if;
        axi_str_txc_tready_int_dly <= axi_str_txc_tready_int;
      end if;
    end process;

    AXI_STR_TXC_TREADY <= axi_str_txc_tready_int;  --fix me  need to look at all txc control and TDX tlast

    -----------------------------------------------------------------------------
    --  Register and hold the axi_flag information and CSUM Control information
    --    axi_flag
    --      0x5 = Status control
    --      0xA = Normal control
    --      0xF = Null Control
    --    CSUM
    --      00 = No CSUM will be performed
    --      01 = Partial Checksum will be performed
    --      10 = Full checksum offloading will be performed
    -----------------------------------------------------------------------------
    CNTRL_WD0 : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          axi_flag   <= (others => '0');
        elsif set_axi_flag = '1' then
          axi_flag   <= axi_str_txc_tdata_dly0(31 downto 28);
        else
          axi_flag   <= axi_flag;
        end if;
      end if;
    end process;

    CNTRL_WD1 : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          csum_cntrl <= (others => '0');
        elsif set_csum_cntrl = '1' then
          csum_cntrl <= axi_str_txc_tdata_dly0 (1 downto  0);
        else
          csum_cntrl <= csum_cntrl;
        end if;
      end if;
    end process;

      ---------------------------------------------------------------------------
      --  Delay signal to load csum value in csum calculation
      ---------------------------------------------------------------------------
      CHECK_FULL_SIG : process(AXI_STR_TXC_ACLK)
      begin

        if rising_edge(AXI_STR_TXC_ACLK) then
          check_full <= set_txc_addr_4_n;
        end if;
      end process;


    -----------------------------------------------------------------------------
    --  This generate is used to reduce a small amount of logic when the CSUM
    --    functionality is not included in the build
    -----------------------------------------------------------------------------
    GEN_CSUM_SUPPORT : if C_TXCSUM /= 0 generate
    begin

      ---------------------------------------------------------------------------
      --  Used when C_CSUM = 1 and the csum_cntrl=01 in the AXI Stream Control
      --    Word 0
      --      csum_begin tells the HW where to start calculating the CSUM
      --      csum_insert tells the HW where to insert the calculated CSUM
      ---------------------------------------------------------------------------
      CNTRL_WD1 : process(AXI_STR_TXC_ACLK)
      begin

        if rising_edge(AXI_STR_TXC_ACLK) then
          if reset2axi_str_txc = '1' then
            csum_begin_int    <= (others => '0');
            csum_begin_bytes  <= (others => '0');
            csum_insert_int   <= (others => '0');
            csum_insert_bytes <= (others => '0');
          elsif set_csum_begin_insert = '1' then
            csum_begin_int    <= std_logic_vector(unsigned(zeroes_csum & axi_str_txc_tdata_dly0(c_TxD_addrb_width  +17 downto 18)) +
                                                  unsigned(zeroes_csum & axi_str_txd_2_mem_addr_int) - 1);
            csum_begin_bytes  <= axi_str_txc_tdata_dly0(17 downto 16);
            csum_insert_int   <= std_logic_vector(unsigned(zeroes_csum & axi_str_txc_tdata_dly0(c_TxD_addrb_width  + 1 downto  2))  +
                                                  unsigned(zeroes_csum & axi_str_txd_2_mem_addr_int));
            csum_insert_bytes <= axi_str_txc_tdata_dly0( 1 downto  0);
          else
            csum_begin_int    <= csum_begin_int;
            csum_begin_bytes  <= csum_begin_bytes;
            csum_insert_int   <= csum_insert_int;
            csum_insert_bytes <= csum_insert_bytes;
          end if;
        end if;
      end process;

      --  Cannot begin or insert at a value larger than the memory so mask off the unused bits:
      --    32K/4 -> 8K   of addressing -> (12:0)
      --    16K/4 -> 4K   of addressing -> (11:0)
      --     8K/4 -> 2K   of addressing -> (10:0)
      --     4K/4 -> 1K   of addressing -> ( 9:0)
      --     2K/4 -> 512M of addressing -> ( 8:0)
      csum_begin  <= csum_begin_int(c_TxD_addrb_width   -1 downto  0);
      csum_insert <= csum_insert_int(c_TxD_addrb_width   -1 downto  0);

      ---------------------------------------------------------------------------
      --  Used when C_CSUM = 1 and the csum_cntrl=01 in the AXI Stream Control
      --    Word 0
      --      csum_init tells the HW what to initialize the CSUM to before
      --        starting the CSUM calculation
      ---------------------------------------------------------------------------
      CNTRL_WD2 : process(AXI_STR_TXC_ACLK)
      begin

        if rising_edge(AXI_STR_TXC_ACLK) then
          if reset2axi_str_txc = '1' then
            csum_init  <= (others => '0');
          elsif set_csum_rsvd_init = '1' then
            csum_init  <= axi_str_txc_tdata_dly0(15 downto  0);
          else
            csum_init  <= csum_init;
          end if;
        end if;
      end process;


      ---------------------------------------------------------------------------
      --  Delay signal to load csum value in csum calculation
      ---------------------------------------------------------------------------
      CSUM_INIT_LOAD : process(AXI_STR_TXC_ACLK)
      begin

        if rising_edge(AXI_STR_TXC_ACLK) then
          if set_csum_rsvd_init = '1' then
            load_csum_int <= '1';
          else
            load_csum_int <= '0';
          end if;
        end if;
      end process;

      csum_addr <= axi_str_txd_2_mem_addr_int;



      I_TX_CSUM : tx_csum_partial_calc_if
      generic map (
        C_FAMILY                  => C_FAMILY,
        C_TXCSUM                  => C_TXCSUM,
        C_S_AXI_DATA_WIDTH        => C_S_AXI_DATA_WIDTH,
        c_TxD_addrb_width         => c_TxD_addrb_width
      )
      port map (
        AXI_STR_TXC_ACLK           => AXI_STR_TXC_ACLK,
        reset2axi_str_txc          => reset2axi_str_txc,
        axi_str_txc_tready_int_dly => axi_str_txc_tready_int_dly,
        axi_str_txc_tvalid_dly0    => axi_str_txc_tvalid_dly0,
        axi_str_txc_tlast_dly0     => axi_str_txc_tlast_dly0,

        load_csum_int              => load_csum_int,
        axi_flag                   => axi_flag,
        csum_cntrl                 => csum_cntrl,
        csum_begin                 => csum_begin,
        csum_begin_bytes           => csum_begin_bytes,
        csum_insert                => csum_insert,
        csum_insert_bytes          => csum_insert_bytes,
        csum_init                  => csum_init,

        AXI_STR_TXD_ACLK           => AXI_STR_TXD_ACLK,
        reset2axi_str_txd          => reset2axi_str_txd,
        csum_addr                  => csum_addr,
        inc_txd_wr_addr            => inc_txd_wr_addr,
        inc_txd_addr_one           => inc_txd_addr_one,
        non_xilinx_ip_pulse        => '0',
        axi_str_txd_tdata_dly1     => axi_str_txd_tdata_dly1,

        do_csum                    => do_csum,
        csum_result                => csum_result,
        csum_en                    => csum_en,
        csum_we                    => csum_we,
        csum_cmplt                 => csum_cmplt
      );


    end generate GEN_CSUM_SUPPORT;


    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Data Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXD_CONTROL : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_tvalid_dly0 <= '0';
          axi_str_txd_tlast_dly0  <= '0';
          clr_txd_trdy            <= '0';
        else
          axi_str_txd_tvalid_dly0 <= AXI_STR_TXD_TVALID;
          axi_str_txd_tlast_dly0  <= AXI_STR_TXD_TLAST;
          if axi_str_txd_tvalid = '1' and axi_str_txd_tlast = '1' and axi_str_txd_tready_int = '1' then
            clr_txd_trdy <= '1';
          else
            clr_txd_trdy <= '0';
          end if;
        end if;
      end if;
    end process;

    AXI_STR_TXD_TREADY <= axi_str_txd_tready_int;  --fix me  need to look at all txd control and TXC tlast

    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Data Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXD_IN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_tstrb_dly0  <= AXI_STR_TXD_TSTRB;
        axi_str_txd_tdata_dly0  <= AXI_STR_TXD_TDATA;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Delay the data one more clock for BRAM
    -----------------------------------------------------------------------------
    REG_TXD_DLY0 : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if csum_en = '1' then
        -- Mux in the CSUM result
        --  The WE will only allow a 16 bit write to memory
          axi_str_txd_tdata_dly1 <= csum_result(15 downto 0) & csum_result(15 downto 0);
        elsif axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
        -- Zero out invalid data so CSUM calculation is correct
          case axi_str_txd_tstrb_dly0 is
            when "0000" => axi_str_txd_tdata_dly1  <= (others => '0');
            when "0001" => axi_str_txd_tdata_dly1  <= X"000000" & axi_str_txd_tdata_dly0( 7 downto 0);
            when "0011" => axi_str_txd_tdata_dly1  <= X"0000"   & axi_str_txd_tdata_dly0(15 downto 0);
            when "0111" => axi_str_txd_tdata_dly1  <= X"00"     & axi_str_txd_tdata_dly0(23 downto 0);
            when others => axi_str_txd_tdata_dly1  <=             axi_str_txd_tdata_dly0;
          end case;
        else
          axi_str_txd_tdata_dly1  <= axi_str_txd_tdata_dly1;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  AXI Stream TX Data State Machine - combinational/combinatorial
    --    Used to provide the control to write the data to the BRAM
    --    This state machine will throttle the Transmit AXI Stream Control state
    --      machine until after the data information has been received.
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXD_CMB : process (txd_wr_cs,axi_str_txd_tvalid_dly0,
      axi_str_txd_tlast_dly0,
      axi_str_txd_tstrb_dly0,wrote_first_packet,axi_str_txd_tready_int_dly,
      txd_rd_pntr,txd_mem_full,txd_min_wr_addr,
      txd_rd_pntr_hold,do_csum,txd_rdy,csum_en,txd_mem_afull,txd_rd_pntr_hold_plus3,
      compare_addr0_cmplt,
      axi_str_txd_2_mem_addr_int,txd_max_wr_addr,
      check_full,txd_max_wr_addr_minus4)
    begin

      inc_txd_wr_addr     <= '0';
      set_txd_we          <= "0000";
      set_txd_en          <= '0';
      set_first_packet    <= '0';
      set_txd_rdy         <= '0';
      clr_txd_rdy         <= '0';
      clr_full_pntr       <= '0';
      disable_txd_trdy    <= '0';
      disable_txc_trdy    <= '0';
      halt_pntr_update    <= '0';
      set_txd_mem_full    <= '0';
      clr_txd_mem_full    <= '0';
      set_txd_mem_afull   <= '0';
      update_rd_pntrs     <= '0';

      case txd_wr_cs is
        when IDLE =>
          if compare_addr0_cmplt = '1' then
          --  Requirement is that the TXD and TXC interfaces use the same clock
          --    so it is OK to used the TXC signals in the TXD state machine
            set_txd_rdy <= '1';
            txd_wr_ns   <= TXD_PRM;
          else
            set_txd_rdy <= '0';
            txd_wr_ns   <= IDLE;
          end if;
        when TXD_PRM =>
--      Made change to ensure TxD Memory is never full here.
--      The memory can always accept data at the start of a transfer
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
          --  delay incrementing pointer until next data
          --    Ethernet has to send 14bytes as a bare minimum, so it is
          --    guaranteed to get through this state with all of the strobes set
          --    and TLAST = '0'
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            disable_txd_trdy    <= '0';
            txd_wr_ns           <= TXD_WRT;
          else
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            disable_txd_trdy    <= '0';
            txd_wr_ns           <= TXD_PRM;
          end if;
        when  TXD_WRT =>
          if txd_mem_full = '1' and axi_str_txd_tready_int_dly = '0' then
          --memory is full when axi_str_txd_tready_int_dly = '0'
            inc_txd_wr_addr     <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_first_packet    <= '0';
            clr_txd_rdy         <= '0';
            disable_txd_trdy    <= '1';
            txd_wr_ns           <= MEM_FULL;
          elsif axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
            inc_txd_wr_addr     <= '1';
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            if axi_str_txd_tlast_dly0 = '1' then
              if do_csum = '1' then
              --  do not care if memory is full because we are over-writing
              --  a location
                set_first_packet    <= '0';
                clr_txd_rdy         <= '1';
                disable_txc_trdy    <= '1';
                disable_txd_trdy    <= '0';
                txd_wr_ns           <= WAIT_CSUM;
              else-- txd_mem_full = '1' or txd_mem_afull = '1'
              --  received TLAST but fifo is full so wait until it can
              --  accept more data before going idle

                if wrote_first_packet = '0' then
                  set_first_packet <= '1';
                else
                  set_first_packet <= '0';
                end if;

                clr_txd_rdy         <= '1';
                disable_txc_trdy    <= '1';
                disable_txd_trdy    <= '0';
                txd_wr_ns           <= WAIT_WR1;
              end if;
            else
            --  received data (normal receive), so continue receiving data
              set_first_packet    <= '0';
              clr_txd_rdy         <= '0';
              disable_txd_trdy    <= '0';
              txd_wr_ns           <= TXD_WRT;
            end if;
          else
            inc_txd_wr_addr     <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_first_packet    <= '0';
            clr_txd_rdy         <= '0';
            disable_txd_trdy    <= '0';
            txd_wr_ns           <= TXD_WRT;
          end if;
       when MEM_FULL =>
          --  stay here until the read pointer updates by 4 words or more.  The read side operates on bytes,
          --  the write side operates on words.
          --    The read pointer updates every 512 bytes (128 words) and at the end of a packet.
          --      The samallest packet the can be sent is 15bytes, but since the BRAM is 32 bit aligned,
          --      the read side will usually update the read pointer by a minimum of 16 bytes (4 words).  However,
          --      it can update by by less than 16 bytes (4 words).  This can occure if a packet started at read
          --      address 0x1A4 (write address 0x69), and the packet is 516 bytes in length (129 words).  Here the read pointer
          --      will update at 0x3A4 (write address 0xE9 - 128 words) then again at the end of the packet at 0x3A8
          --      (write address 0xEA).
          --        If this occures the below logic will detect it and update the read pointer, but stay in this
          --        state until the next update occurs.  The next update is guaranteed to be greater than 4 words,
          --        which will allow the full pointers to be cleared for the next packet.
          inc_txd_wr_addr     <= '0';
          set_txd_we          <= "0000";
          set_txd_en          <= '0';
          set_first_packet    <= '0';
          clr_txd_rdy         <= '0';
          if txd_rd_pntr = txd_rd_pntr_hold then
          --  stay here until an update occurs
            update_rd_pntrs  <= '0';
            disable_txd_trdy <= '1';
            clr_full_pntr    <= '0';
            txd_wr_ns        <= MEM_FULL;
          else
          --  The read pointer was updated to determine if it was updated by 4 words or more
          --    If not, update the hold pointers, but stay in this state
            if txd_rd_pntr_hold <= txd_max_wr_addr_minus4 then
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x0 - 0x1FB
              if txd_rd_pntr > txd_rd_pntr_hold_plus3 then
              -- an update of 4 words or greater occured so exit this state
                update_rd_pntrs  <= '0';
                disable_txd_trdy <= '0';
                clr_full_pntr    <= '1';
                txd_wr_ns        <= TXD_WRT;
              else
              --  the update was less than 4 words
              --    (txd_rd_pntr <= txd_rd_pntr_hold_plus3)
                if txd_rd_pntr < txd_rd_pntr_hold then
                --  the read pointer wrapped, so exit because the update was > 4 words
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              end if;
            else
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x1FC- 0x1FF
              if txd_rd_pntr_hold_plus3 = txd_max_wr_addr then
              --  txd_rd_pntr = 0x1FC for 2048 byte memory, so txd_rd_pntr_hold_plus3 = max memory size
                if (txd_rd_pntr <= txd_rd_pntr_hold) then
                --  the update was >= 4 words so exit
                --    for a 2048 memory, txd_rd_pntr_hold = 0x1FC
                --      if txd_rd_pntr is between 0x0 and 0x1FB then an update of 4 or more words occurred
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              else
              --  txd_rd_pntr = 0x1FD, 0x1FE, or 0x1FF for 2048 byte memory,
              --  so the minimum txd_rd_pntr_hold_plus3 can be is 0, 1, or 2
                if (txd_rd_pntr > txd_rd_pntr_hold_plus3) and (txd_rd_pntr < txd_rd_pntr_hold) then
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr has to be tween 0x1 and 0x1FC to exit this state
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr has to be tween 0x2 and 0x1FD to exit this state
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr has to be tween 0x3 and 0x1FE to exit this state
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  txd_rd_pntr did not update by 4 or more words, so update hold poointers and stay in this state
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited BUT
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr was only updated 1-3 words to 0x1FE, 0x1FF, or 0x0, so stay here
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr was only updated 1-3 words to 0x1FF, 0x0, or 0x1, so stay here
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr was only updated 1-3 words to 0x0, 0x1, or 0x2, so stay here
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              end if;
            end if;
          end if;

        when CLR_FULL =>
          --  stay here until the read pointer updates by 4 words or more.  The read side operates on bytes,
          --  the write side operates on words.
          --    The read pointer updates every 512 bytes (128 words) and at the end of a packet.
          --      The samallest packet the can be sent is 15bytes, but since the BRAM is 32 bit aligned,
          --      the read side will usually update the read pointer by a minimum of 16 bytes (4 words).  However,
          --      it can update by by less than 16 bytes (4 words).  This can occure if a packet started at read
          --      address 0x1A4 (write address 0x69), and the packet is 516 bytes in length (129 words).  Here the read pointer
          --      will update at 0x3A4 (write address 0xE9 - 128 words) then again at the end of the packet at 0x3A8
          --      (write address 0xEA).
          --        If this occures the below logic will detect it and update the read pointer, but stay in this
          --        state until the next update occurs.  The next update is guaranteed to be greater than 4 words,
          --        which will allow the full pointers to be cleared for the next packet.
          inc_txd_wr_addr     <= '0';
          set_txd_we          <= "0000";
          set_txd_en          <= '0';
          set_first_packet    <= '0';
          clr_txd_rdy         <= '0';
          if txd_rd_pntr = txd_rd_pntr_hold then
          --  stay here until an update occurs
            update_rd_pntrs  <= '0';
            halt_pntr_update <= '1';
            disable_txc_trdy <= '1';
            disable_txd_trdy <= '1';
            clr_full_pntr    <= '0';
            txd_wr_ns        <= CLR_FULL;
          else
          --  The read pointer was updated to determine if it was updated by 4 words or more
          --    If not, update the hold pointers, but stay in this state
            if txd_rd_pntr_hold <= txd_max_wr_addr_minus4 then
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x0 - 0x1FB
              if txd_rd_pntr > txd_rd_pntr_hold_plus3 then
              -- an update of 4 words or greater occured so exit this state
                if wrote_first_packet = '0' then
                  set_first_packet <= '1';
                else
                  set_first_packet <= '0';
                end if;
                update_rd_pntrs  <= '0';
                halt_pntr_update <= '0';
                disable_txd_trdy <= '0';
                clr_full_pntr    <= '1';
                clr_txd_rdy      <= '0';
                txd_wr_ns        <= WAIT_COMPARE_CMPLT;
              else
              --  the update was less than 4 words
              --    (txd_rd_pntr <= txd_rd_pntr_hold_plus3)
                if txd_rd_pntr < txd_rd_pntr_hold then
                --  the read pointer wrapped, so exit because the update was > 4 words
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  halt_pntr_update <= '1';
                  disable_txc_trdy <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= CLR_FULL;
                end if;
              end if;
            else
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x1FC- 0x1FF
              if txd_rd_pntr_hold_plus3 = txd_max_wr_addr then
              --  txd_rd_pntr = 0x1FC for 2048 byte memory, so txd_rd_pntr_hold_plus3 = max memory size
                if (txd_rd_pntr <= txd_rd_pntr_hold) then
                --  the update was >= 4 words so exit
                --    for a 2048 memory, txd_rd_pntr_hold = 0x1FC
                --      if txd_rd_pntr is between 0x0 and 0x1FB then an update of 4 or more words occurred
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  halt_pntr_update <= '1';
                  disable_txc_trdy <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= CLR_FULL;
                end if;
              else
              --  txd_rd_pntr = 0x1FD, 0x1FE, or 0x1FF for 2048 byte memory,
              --  so the minimum txd_rd_pntr_hold_plus3 can be is 0, 1, or 2
                if (txd_rd_pntr > txd_rd_pntr_hold_plus3) and (txd_rd_pntr < txd_rd_pntr_hold) then
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr has to be tween 0x1 and 0x1FC to exit this state
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr has to be tween 0x2 and 0x1FD to exit this state
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr has to be tween 0x3 and 0x1FE to exit this state
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  txd_rd_pntr did not update by 4 or more words, so update hold poointers and stay in this state
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited BUT
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr was only updated 1-3 words to 0x1FE, 0x1FF, or 0x0, so stay here
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr was only updated 1-3 words to 0x1FF, 0x0, or 0x1, so stay here
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr was only updated 1-3 words to 0x0, 0x1, or 0x2, so stay here
                  update_rd_pntrs  <= '1';
                  halt_pntr_update <= '1';
                  disable_txc_trdy <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= CLR_FULL;
                end if;
              end if;
            end if;
          end if;

        when WAIT_CSUM =>
          if txd_mem_full = '1' then -- hold until complete with CSUM
            set_txd_mem_full <= '1';
          else
            set_txd_mem_full <= '0';
          end if;

          if txd_mem_afull = '1' then -- hold until complete with CSUM
            set_txd_mem_afull <= '1';
          else
            set_txd_mem_afull <= '0';
          end if;

          if csum_en = '1' then --one clock cycle pulse - asserts on 4th clock cycle in this state
            if txd_mem_full = '1' or txd_mem_afull = '1' then
              set_first_packet  <= '0';
              disable_txc_trdy  <= '1';
              disable_txd_trdy  <= '1';
              clr_txd_mem_full  <= '0';
              txd_wr_ns         <= CLR_FULL;
            else
              if wrote_first_packet = '0' then
                set_first_packet <= '1';
              else
                set_first_packet <= '0';
              end if;
              set_first_packet  <= '0';
              disable_txc_trdy  <= '0';
              disable_txd_trdy  <= '0';
              clr_txd_mem_full  <= '0';
              txd_wr_ns         <= IDLE;
            end if;
          else
            clr_txd_rdy       <= '0';
            disable_txc_trdy  <= '1';
            clr_txd_mem_full  <= '0';
            txd_wr_ns         <= WAIT_CSUM;
          end if;

        when WAIT_WR1 =>
          disable_txc_trdy  <= '1';
          disable_txd_trdy  <= '0';

          if check_full = '1' then
            txd_wr_ns         <= WAIT_WR2;
          else
            txd_wr_ns         <= WAIT_WR1;
          end if;
        when WAIT_WR2 =>
          if txd_mem_full = '1' or txd_mem_afull = '1' then
            disable_txc_trdy  <= '1';
            disable_txd_trdy  <= '1';
            txd_wr_ns         <= CLR_FULL;
          else
            if wrote_first_packet = '0' then
              set_first_packet <= '1';
            else
              set_first_packet <= '0';
            end if;

            disable_txc_trdy  <= '0';
            disable_txd_trdy  <= '0';
            txd_wr_ns         <= IDLE;
          end if;
        when WAIT_COMPARE_CMPLT =>
          txd_wr_ns        <= IDLE;
        when others =>
          txd_wr_ns <= IDLE;
      end case;
    end process;

    -----------------------------------------------------------------------------
    -- AXI Stream TX Control State Machine Sequencer
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXD_SEQ : process (AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_wr_cs <= IDLE;
        else
          txd_wr_cs <= txd_wr_ns;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    -- Indicator when performing a write to TxD Memory
    --  clear on axi_str_txd_tlast_dly0 = '1'
    -----------------------------------------------------------------------------
    TXD_RDY_INDICATOR : process (AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rdy <= '0';
        else
          if clr_txd_rdy = '1' then
            txd_rdy <= '0';
          elsif set_txd_rdy = '1' then
            txd_rdy <= '1';
          else
            txd_rdy <= txd_rdy;
          end if;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Filter to indicate first packet was written
    --    Needed for full flag
    -----------------------------------------------------------------------------
    FIRST_PACKET_WROTE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          wrote_first_packet <= '0';
        elsif set_first_packet = '1' then
          wrote_first_packet <= '1';
        else
          wrote_first_packet <= wrote_first_packet;
        end if;
      end if;
    end process;


    axi_str_txd_2_mem_addr_int_plus1 <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 1);
    axi_str_txd_2_mem_addr_int_plus2 <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 2);
    axi_str_txd_2_mem_addr_int_plus3 <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 3);
    axi_str_txd_2_mem_addr_int_plus4 <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 4);


    ---------------------------------------------------------------------------
    --  Register to help fmax
    --  With ASYNC BRAM clock cannot read/write same address in memory at same
    --  time unless timing is met, so read until data matches
    ---------------------------------------------------------------------------
    RD_PNTR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rd_pntr_1 <= (others => '0');
          txd_rd_pntr   <= (others => '0');
          compare_addr0_cmplt <= '0';
        else
          if set_txc_addr_0 = '1' and txc_addr_0_dly2 = '1' and
             txc_we_dly2 = '0'  then
          --  txc_addr_0_dly2 is when data is first avaliable from memory

          --  use set_txc_addr_0 to disable compare_addr0_cmplt once pointers update
          --  once state machine advances, set_txc_addr_0 will go low so use it to disable any more
          --  any more data from memory
            txd_rd_pntr_1      <= Axi_Str_TxC_2_Mem_Dout(c_TxD_addrb_width -1 downto 0);

            if Axi_Str_TxC_2_Mem_Dout(c_TxD_addrb_width -1 downto 0) = txd_rd_pntr_1 and
              compare_addr0_cmplt = '0' then
              txd_rd_pntr         <= txd_rd_pntr_1;
              if enable_compare_addr0_cmplt = '1' then
                compare_addr0_cmplt <= '1';
              else
                compare_addr0_cmplt <= '0';
              end if;
            else
              txd_rd_pntr         <= txd_rd_pntr;
              compare_addr0_cmplt <= '0';
            end if;
          else
            txd_rd_pntr_1      <= txd_rd_pntr_1;
            txd_rd_pntr        <= txd_rd_pntr;
            compare_addr0_cmplt<= '0';
          end if;
        end if;
      end if;
    end process;


    ---------------------------------------------------------------------------
    --  Update the read pointer locations until the memory goes FULL
    --    Then use the stored values to compare against real time read pointer
    --    and throttle appropriately
    ---------------------------------------------------------------------------
    RD_PNTRS : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rd_pntr_hold_plus3 <= txc_rd_addr3;
          txd_rd_pntr_hold       <= txc_rd_addr0;
        else
          if (txd_mem_full = '0' and txc_addr_0_dly2 = '1' and halt_pntr_update = '0') or update_rd_pntrs = '1'then -- wait on this as it might not be needed  or update_hold_pntrs = '1' then --and
          --  halt_pntr_update is for the special case when memory is almost full/full and
          --  the Txd FSM needs to wait for a few reads before the next packet starts
          --  The TxD FSM will assert it HIGH to prevent the poiners from being updated
            txd_rd_pntr_hold_plus3 <= std_logic_vector(unsigned(txd_rd_pntr) +3);
            txd_rd_pntr_hold       <= txd_rd_pntr;
          else
            txd_rd_pntr_hold_plus3 <= txd_rd_pntr_hold_plus3;
            txd_rd_pntr_hold       <= txd_rd_pntr_hold;
          end if;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Full flag indicator
    --    Does not begin comparison until 1st packet is written to memory
    -----------------------------------------------------------------------------
    TXD_FULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
            txd_mem_full     <= '0';
            txd_mem_not_full <= '1';
        else
            if (axi_str_txd_2_mem_addr_int_plus3 = txd_rd_pntr and
                (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) or
               set_txd_mem_full = '1' then
              txd_mem_full     <= '1';
              txd_mem_not_full <= '0';
            else
              txd_mem_full     <= txd_mem_full;
              txd_mem_not_full <= txd_mem_not_full;
            end if;
        end if;
      end if;
    end process;

    TXD_AFULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
            txd_mem_afull     <= '0';
        else

          if (axi_str_txd_2_mem_addr_int_plus4 = txd_rd_pntr and
              (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) or
             set_txd_mem_afull = '1' then
            txd_mem_afull     <= '1';
          else
            txd_mem_afull     <= txd_mem_afull;
          end if;
        end if;
      end if;
    end process;

    DELAY_TXD_TREADY_DISABLE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        disable_txd_trdy_dly <= disable_txd_trdy;
      end if;
    end process;

    DELAY_TREADY_DISABLE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        disable_txc_trdy_dly <= disable_txc_trdy;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  TxD Ready
    --    Only assert when FIFO is not full and TxC is not in process
    -----------------------------------------------------------------------------
    TXD_READY : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_tready_int_dly <= axi_str_txd_tready_int;
        if (AXI_STR_TXD_TLAST = '1' and AXI_STR_TXD_TVALID = '1' and axi_str_txd_tready_int = '1') or
           (clr_txd_trdy = '1' and disable_txd_trdy_dly = '0') or
           disable_txd_trdy = '1' then
          axi_str_txd_tready_int <= '0';
        elsif set_txd_rdy = '1' or (txd_rdy = '1' and clr_txd_rdy = '0') then
            if (axi_str_txd_2_mem_addr_int_plus3 = txd_rd_pntr and
               inc_txd_wr_addr = '1') or
               (clr_full_pntr = '0' and txd_mem_full = '1') then
            --  txd_rd_pntr is where the the current read is occuring, so
            --    to account for register pipelines, this needs to stop at
            --    3 counts before the current write address
              axi_str_txd_tready_int <= '0';
            else
              axi_str_txd_tready_int <= '1';
            end if;
        else
          axi_str_txd_tready_int <= '0';
        end if;
      end if;
    end process;

    AXI_STR_TXD_TREADY     <= axi_str_txd_tready_int;


    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_WR_ADDR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_2_mem_addr_int       <= (others => '0');
          axi_str_txd_2_mem_addr_int_mins1 <= (others => '0');
        elsif (inc_txd_wr_addr = '1' or inc_txd_addr_one = '1') then
        --  the address ready for the next transaction
          axi_str_txd_2_mem_addr_int       <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 1);
          axi_str_txd_2_mem_addr_int_mins1 <= axi_str_txd_2_mem_addr_int;
        elsif csum_en = '1' then
          axi_str_txd_2_mem_addr_int       <= csum_insert(c_TxD_addrb_width   -1 downto 0);
          axi_str_txd_2_mem_addr_int_mins1 <= axi_str_txd_2_mem_addr_int_mins1;
        elsif csum_en_dly = '1' then
          axi_str_txd_2_mem_addr_int       <= axi_str_txd_2_mem_addr_int_last;
          axi_str_txd_2_mem_addr_int_mins1 <= axi_str_txd_2_mem_addr_int_mins1;
        else
          axi_str_txd_2_mem_addr_int       <= axi_str_txd_2_mem_addr_int;
          axi_str_txd_2_mem_addr_int_mins1 <= axi_str_txd_2_mem_addr_int_mins1;
        end if;
      end if;
    end process;


    ---------------------------------------------------------------------------
    --  Force and update the BRAM with the axi_str_txd_2_mem_addr_int
    --  every ~128 writes (~512 bytes)
    ---------------------------------------------------------------------------
    BRAM_UPDATE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_txd_rdy = '1' then
          update_bram_cnt     <= (others => '0');
        else
          if update_bram_cnt(7) = '1' and inc_txd_wr_addr = '1' then
            update_bram_cnt <= unsigned('0' & update_bram_cnt(6 downto 0)) + 1;
          elsif inc_txd_wr_addr = '1' then
            update_bram_cnt <= update_bram_cnt + 1;
          else
            update_bram_cnt <= update_bram_cnt;
          end if;
        end if;
      end if;
    end process;



    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_WR_ADDR_LAST : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_2_mem_addr_int_last <= (others => '0');
        elsif csum_en = '1' then
        --  hold TxD address to restore after CSUM is written
          axi_str_txd_2_mem_addr_int_last <= axi_str_txd_2_mem_addr_int;
        else
          axi_str_txd_2_mem_addr_int_last <= axi_str_txd_2_mem_addr_int_last;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay the CSUM enable to resore the memory address after the CSUM value
    --  is written
    -----------------------------------------------------------------------------
    CSUM_ENABLE_DELAY : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        csum_en_dly <= csum_en;
      end if;
    end process;


    axi_str_txd_2_mem_addr               <= axi_str_txd_2_mem_addr_int;


    Axi_Str_TxD_2_Mem_Din(35)           <= axi_str_txd_2_mem_we_int(3);
    Axi_Str_TxD_2_Mem_Din(26)           <= axi_str_txd_2_mem_we_int(2);
    Axi_Str_TxD_2_Mem_Din(17)           <= axi_str_txd_2_mem_we_int(1);
    Axi_Str_TxD_2_Mem_Din(8)            <= axi_str_txd_2_mem_we_int(0);

    Axi_Str_TxD_2_Mem_Din(34 downto 27) <= axi_str_txd_tdata_dly1(31 downto 24);
    Axi_Str_TxD_2_Mem_Din(25 downto 18) <= axi_str_txd_tdata_dly1(23 downto 16);
    Axi_Str_TxD_2_Mem_Din(16 downto  9) <= axi_str_txd_tdata_dly1(15 downto  8);
    Axi_Str_TxD_2_Mem_Din(7  downto  0) <= axi_str_txd_tdata_dly1( 7 downto  0);

    -----------------------------------------------------------------------------
    --  Write Parity bits to the AXI Stream Data Memory
    --    The parity bit always should be the AXI_STR_TXD_TSTRB bits delayed
    --    except when writing the CSUM value.  If writing CSUM, these bits need
    --    set HIGH for the Half word being written; otherwise, the transmission
    --    will end prematurely.
    -----------------------------------------------------------------------------
    MEM_TXD_PARITY : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if csum_en = '1' then
          axi_str_txd_2_mem_we_int <= csum_we;
        else
          axi_str_txd_2_mem_we_int <= set_txd_we;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Write Enable bits to the AXI Stream Data Memory
    --    All of the write enables bits should be forced HIGH any time a write to
    --    memory is being performed (except csum).  This will allow the parity
    --    bits to be cleared which in turn prevents too much data being read on
    --    the Txd client interface.
    --  When CSUM is being performed, only set the WEs for the half word being
    --  accessed.
    -----------------------------------------------------------------------------
    MEM_TXD_WR_EN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if csum_en = '1' then
          Axi_Str_TxD_2_Mem_We <= csum_we;
        else
          case set_txd_we is
            when "0000" => Axi_Str_TxD_2_Mem_We <= "0000";
            when others => Axi_Str_TxD_2_Mem_We <= "1111";
          end case;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Enable bit to the AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_EN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if set_txd_en = '1' or csum_en = '1' then
          axi_str_txd_2_mem_en_int <= '1';
        else
          axi_str_txd_2_mem_en_int <= '0';
        end if;
      end if;
    end process;

    Axi_Str_TxD_2_Mem_En <= axi_str_txd_2_mem_en_int;

-------------------------------------------------------------------------------
--  End Partial CSUM
-------------------------------------------------------------------------------

end rtl;


-------------------------------------------------------------------------------
-- tx_csum_full_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_csum_full_if.vhd
-- Version:         v1.00a
-- Description:     embedded ip AXI Stream transmit interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--                    tx_axistream_if.vhd
--                      tx_basic_if.vhd
--                      tx_csum_if.vhd
--          ->            tx_csum_full_if.vhd
--                          tx_csum_full_fsm.vhd
--                          tx_csum_full_calc_if.vhd
--                        tx_partial_csum_if.vhd
--                          tx_csum_partial_calc_if.vhd
--                      tx_vlan_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tx_if_pack.all;

-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity tx_csum_full_if is
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data


    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0)   --  Tx AXI-Stream Control to Memory Full Flag

  );

end tx_csum_full_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of tx_csum_full_if is


-------------------------------------------------------------------------------
--  Start Full CSUM
-------------------------------------------------------------------------------
  constant zeroes_txc                     : std_logic_vector(c_TxC_write_width_b -1 downto c_TxC_addrb_width) := (others => '0');
  constant zeroes_txd                     : std_logic_vector(c_TxC_write_width_b -1 downto c_TxD_addrb_width) := (others => '0');
  constant zeroes_txd_2                   : std_logic_vector(c_TxC_write_width_b -1 downto c_TxD_addrb_width + 2 ) := (others => '0');

  type TXC_WR_FSM_TYPE is (
                       TXC_ADDR2_WR,
                       TXC_ADDR0_WR,
                       WAIT_WR_CMPLT,
                       TXC_WD0,
--                       WAIT_TXD_FULL,
                       TXC_WD1,
                       WAIT_ADDR2_COMPARE_CMPLT,--added for BRAM async clocks
                       TXC_WD2,
                       TXC_WD3,
                       TXC_WD4,
                       WAIT_ADDR0_COMPARE_CMPLT,--added for BRAM async clocks
                       TXC_WD5,
                       WAIT_TXD_CMPLT,
                       WAIT_TXD_MEM,
                       WR_TXC_PNTR,
                       WAIT_CSUM_END,
                       WR_TXD_END_PNTR
                      );
  signal txc_wr_cs, txc_wr_ns             : TXC_WR_FSM_TYPE;

  type TXD_WR_FSM_TYPE is (
                       IDLE,
                       TXD_PRM,
                       TXD_WRT,
                       MEM_FULL,
                       CLR_FULL,
                       WAIT_WR1,
                       WAIT_WR2,
                       WAIT_CSUM,
                       WAIT_COMPARE_CMPLT
                      );
  signal txd_wr_cs, txd_wr_ns             : TXD_WR_FSM_TYPE;

  signal txc_min_wr_addr                  : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_rsvd_wr_addr                 : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_max_wr_addr                  : std_logic_vector(c_TxC_addrb_width -1 downto 0);

  signal txc_wr_addr0                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr1                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr2                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr3                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr5                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr6                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);

  signal axi_str_txc_tready_int           : std_logic;
  signal axi_str_txc_tready_int_dly       : std_logic;
  signal axi_str_txc_tvalid_dly0          : std_logic;
  signal axi_str_txc_tlast_dly0           : std_logic;
--  signal axi_str_txc_tstrb_dly0           : std_logic_vector(3 downto 0);
  signal axi_str_txc_tdata_dly0           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal clr_txc_trdy                     : std_logic;

  signal axi_str_txd_tready_int           : std_logic;
  signal axi_str_txd_tready_int_dly       : std_logic;
  signal axi_str_txd_tvalid_dly0          : std_logic;
  signal axi_str_txd_tlast_dly0           : std_logic;
  signal axi_str_txd_tstrb_dly0           : std_logic_vector(3 downto 0);
  signal axi_str_txd_tdata_dly0           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal axi_str_txd_tdata_dly1           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal clr_txd_trdy                     : std_logic;

  signal set_txc_addr_0                   : std_logic;
  signal txc_addr_0_dly1                  : std_logic;
  signal txc_addr_0_dly2                  : std_logic;
  signal set_txc_addr_1                   : std_logic;
  signal txc_addr_1                       : std_logic;
  signal set_txc_addr_2                   : std_logic;
  signal txc_addr_2                       : std_logic;
  signal set_txc_addr_4_n                 : std_logic;
  signal set_txc_addr_3                   : std_logic;
  signal clr_txc_addr_3                   : std_logic;
  signal txc_addr_3_dly                   : std_logic;
  signal txc_addr_3_dly2                  : std_logic;
  signal txc_addr_3_dly3                  : std_logic;
  signal inc_txd_addr_one                 : std_logic;
  signal set_txc_trdy                     : std_logic;
  signal set_txc_trdy2                    : std_logic;
  signal clr_txc_trdy2                    : std_logic;
  signal set_txcwr_rd_addr                : std_logic;
  signal set_txcwr_wr_end                 : std_logic;
  signal set_txc_en                       : std_logic;
  signal set_txc_we                       : std_logic;
  signal txc_we                           : std_logic;
  signal txc_we_dly1                      : std_logic;
  signal txc_we_dly2                      : std_logic;

  signal addr_2_en                        : std_logic;
  signal addr_2_en_dly1                   : std_logic;
  signal addr_2_en_dly2                   : std_logic;

  signal txc_mem_full                     : std_logic;
  signal txc_mem_not_full                 : std_logic;
  signal txc_mem_afull                    : std_logic;
  signal txc_mem_wr_addr                  : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_0                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_1                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_last             : std_logic_vector(c_TxC_addrb_width   -1 downto 0);

  signal Axi_Str_TxC_2_Mem_Addr_int       : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal Axi_Str_TxC_2_Mem_We_int         : std_logic_vector(0 downto 0);
  signal txc_mem_wr_addr_plus1            : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_plus2            : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_rd_addr2_pntr                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_rd_addr2_pntr_1              : std_logic_vector(c_TxC_addrb_width   -1 downto 0);


  -- Set to the full width of the write data bus
  signal Axi_Str_TxC_2_Mem_Din_int        : std_logic_vector(c_TxC_write_width_b -1 downto 0);

  signal set_axi_flag                     : std_logic;
  signal set_csum_cntrl                   : std_logic;
  signal set_csum_begin_insert            : std_logic;
  signal set_csum_rsvd_init               : std_logic;
  signal axi_flag                         : std_logic_vector( 3 downto 0);
  signal csum_cntrl                       : std_logic_vector( 1 downto 0);

  signal set_first_packet                 : std_logic;
  signal wrote_first_packet               : std_logic;
  signal inc_txd_wr_addr                  : std_logic;
  signal set_txd_we                       : std_logic_vector( 3 downto 0);
  signal set_txd_en                       : std_logic;
  signal set_txd_rdy                      : std_logic;
  signal clr_txd_rdy                      : std_logic;
  signal clr_full_pntr                    : std_logic;
  signal halt_pntr_update                 : std_logic;
  signal disable_txd_trdy                 : std_logic;
  signal disable_txd_trdy_dly             : std_logic;
  signal disable_txc_trdy                 : std_logic;
  signal disable_txc_trdy_dly             : std_logic;

  signal txd_rdy                          : std_logic;
  signal axi_str_txd_2_mem_addr_int       : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_last  : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_mins1 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus1 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus2 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus3 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus4 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txd_mem_full                     : std_logic;
  signal txd_mem_not_full                 : std_logic;
  signal txd_mem_afull                    : std_logic;
  signal axi_str_txd_2_mem_we_int         : std_logic_vector( 3 downto 0);
  signal axi_str_txd_2_mem_en_int         : std_logic;

  signal txd_rd_pntr                      : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_1                    : std_logic_vector(c_TxD_addrb_width -1 downto 0);

  signal txd_min_wr_addr                  : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_max_wr_addr                  : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_max_wr_addr_minus4           : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_hold_plus3           : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_hold                 : std_logic_vector(c_TxD_addrb_width -1 downto 0);


  signal do_csum                          : std_logic;
--  signal csum_result                      : std_logic_vector(15 downto 0);
  signal csum_en                          : std_logic;
  signal csum_we                          : std_logic_vector(3 downto 0);

  signal csum_en_dly                      : std_logic;
  signal csum_cmplt                       : std_logic;

  signal tx_init_in_prog_int              : std_logic;
  signal init_bram                        : std_logic;

  signal txc_rd_addr0                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txc_rd_addr2                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txc_rd_addr3                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);

  signal set_txd_mem_full                 : std_logic;
  signal clr_txd_mem_full                 : std_logic;
  signal set_txd_mem_afull                : std_logic;

  signal compare_addr0                    : std_logic;
  signal compare_addr0_cmplt              : std_logic;

  signal compare_addr2                    : std_logic;
  signal compare_addr2_cmplt              : std_logic;
  signal compare_addr2_cmplt_dly          : std_logic;

  signal update_bram_cnt                  : unsigned(7 downto 0);

  signal enable_compare_addr0_cmplt       : std_logic;

  --  Full CSUM Signals
  signal abort_csum                       : std_logic;
  signal csum_calc_en                     : std_logic;
  signal clr_csums                        : std_logic;
  signal tcp_ptcl                         : std_logic;
  signal udp_ptcl                         : std_logic;
  signal en_ipv4_hdr_b32                  : std_logic_vector( 1 downto 0);
  signal en_ipv4_hdr_b10                  : std_logic_vector( 1 downto 0);
  signal last_ipv4_hdr_cnt                : std_logic;
  signal hdr_csum_dout                    : std_logic_vector(15 downto 0);  --hook me up
  signal hdr_csum_we                      : std_logic_vector( 3 downto 0);  --hook me up
  signal hdr_csum_cmplt                   : std_logic;                      --hook me up
  signal fsm_csum_en_b32                  : std_logic_vector( 1 downto 0);
  signal fsm_csum_en_b10                  : std_logic_vector( 1 downto 0);
  signal add_psdo_wd                      : std_logic;
  signal ptcl_csum_dout                   : std_logic_vector(15 downto 0);  --hook me up
  signal ptcl_csum_we                     : std_logic_vector( 3 downto 0);  --hook me up
  signal ptcl_csum_cmplt                  : std_logic;                      --hook me up
  signal zeroes_en                        : std_logic_vector( 1 downto 0);
  signal csum_din                         : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal do_ipv4hdr                       : std_logic;
  signal not_tcp_udp                      : std_logic;
  signal do_full_csum                     : std_logic;
  signal wr_hdr_csum                      : std_logic;
  signal wr_ptcl_csum                     : std_logic;
  signal csum_strt_addr                   : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal csum_ipv4_hdr_addr               : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal csum_ipv4_hdr_we                 : std_logic_vector( 3 downto 0);
  signal csum_ptcl_addr                   : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal csum_ptcl_we                     : std_logic_vector( 3 downto 0);
  signal fcsum_fsm_rst                    : std_logic;

  signal inc_txd_addr_one_early           : std_logic;
  signal end_addr_byte_offset             : std_logic_vector(1 downto 0);


  signal check_full                       : std_logic;
  signal update_rd_pntrs                  : std_logic;


  begin

    -----------------------------------------------------------------------------
    --  The TxC BRAM is set up to to always store the current TxD Read and Write
    --    pointers in the first two locations (0x0 and 0x1) of the Memory
    --    respectivively.  The current TxC Read and write pointer are always
    --    stored in the the next two locations (0x2 and 0x3) of the Memory
    --    respectively.  The End addresses for each packet are then stored
    --    in the remaing Memory locations starting at address 0x4.  After
    --    the end pointer to the maximum address has been written, if the
    --    memory is not full, the address pointer will loop back to address
    --    0x4 and write the end pointer for the next packet.
    --
    --                                   BRAM
    --                             Write       Read
    --                           _____________________
    --                          |__________|_________| <-- TxD Rd Pointer
    --      TxD Wr Pointer -->  |__________|_________|
    --                          |__________|_________| <-- TxC Rd Pointer
    --      TxC Wr Pointer -->  |__________|_________|
    --      Packet 0 End   -->  |__________|_________|  --> Packet 0 End
    --      Packet 1 End   -->  |__________|_________|  --> Packet 1 End
    --      Packet 2 End   -->  |__________|_________|  --> Packet 2 End
    --         .                |__________|_________|         .
    --         .                |__________|_________|         .
    --         .                |__________|_________|         .
    --      Packet n End   -->  |__________|_________|  --> Packet n End
    --
    -----------------------------------------------------------------------------

    -----------------------------------------------------------------------------
    --  Create the full and empty comparison values for the S6 and V6 since
    --  1 S6 BRAM = 1/2 V6 BRAM
    -----------------------------------------------------------------------------
    GEN_TXC_MIN_MAX_WR_FLAG : for i in (c_TxC_addrb_width-1) downto 0 generate
      txc_min_wr_addr(i)  <= '1' when (i = 2)          else '0'; -- do not loop back to 0x0; loop to 0x4
      txc_max_wr_addr(i)  <= '0' when (i = 0 or i = 1) else '1';
      txc_wr_addr0(i)     <= '0';
      txc_wr_addr1(i)     <= '1' when (i = 0)          else '0';
      txc_wr_addr2(i)     <= '1' when (i = 1)          else '0';
      txc_wr_addr3(i)     <= '1' when (i = 0 or i = 1) else '0';
      txc_wr_addr5(i)     <= '1' when (i = 0 or i = 2) else '0';
      txc_wr_addr6(i)     <= '1' when (i = 1 or i = 2) else '0';
    end generate GEN_TXC_MIN_MAX_WR_FLAG;

    GEN_TXD_MIN_MAX_WR_FLAG : for i in (c_TxD_addrb_width-1) downto 0 generate
      txd_min_wr_addr(i)        <= '1' when (i = 0) else '0';
      txd_max_wr_addr_minus4(i) <= '0' when (i = 2) else '1';
      txd_max_wr_addr(i)        <= '1';
    end generate GEN_TXD_MIN_MAX_WR_FLAG;


    GEN_TXC_MIN_MAX_RD_FLAG : for i in (c_TxD_addrb_width-1) downto 0 generate
      txc_rd_addr0(i)     <= '0';
      txc_rd_addr2(i)     <= '1' when (i = 1)          else '0';
      txc_rd_addr3(i)     <= '1' when (i = 0 or i = 1) else '0';
    end generate GEN_TXC_MIN_MAX_RD_FLAG;




    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Control Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXC_CONTROL : process(AXI_STR_TXC_ACLK)
    begin
      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          axi_str_txc_tvalid_dly0 <= '0';
          axi_str_txc_tlast_dly0  <= '0';
          clr_txc_trdy           <= '0';
        else
          axi_str_txc_tvalid_dly0 <= axi_str_txc_tvalid;
          axi_str_txc_tlast_dly0  <= axi_str_txc_tlast;
          if axi_str_txc_tvalid = '1' and axi_str_txc_tlast = '1' and axi_str_txc_tready_int = '1' then
            clr_txc_trdy <= '1';
          else
            clr_txc_trdy <= '0';
          end if;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Control Data Bus
    -----------------------------------------------------------------------------
    REG_TXC_IN : process(AXI_STR_TXC_ACLK)
    begin
      if rising_edge(AXI_STR_TXC_ACLK) then
--          axi_str_txc_tstrb_dly0  <= axi_str_txc_tstrb;
          axi_str_txc_tdata_dly0  <= axi_str_txc_tdata;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  AXI Stream TX Control State Machine - combinational/combinatorial
    --    Used to register the incoming control and checksum information
    --    This state machine will throttle the Transmit AXI Stream Data state
    --      machine until after the control information has been received.
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXC_CMB : process (txc_wr_cs,axi_str_txc_tvalid_dly0,
      axi_str_txc_tlast_dly0,axi_str_txd_tlast_dly0,
      axi_str_txd_tvalid_dly0,txc_addr_3_dly,
      wrote_first_packet,axi_str_txc_tready_int_dly,axi_str_txd_tready_int_dly,
      disable_txd_trdy_dly,disable_txc_trdy_dly,do_csum,ptcl_csum_cmplt,
      compare_addr2_cmplt,compare_addr2_cmplt_dly,compare_addr0_cmplt,
      update_bram_cnt,txc_mem_full,
      do_ipv4hdr,do_full_csum)
    begin


      set_axi_flag           <= '0';
      set_csum_cntrl         <= '0';
      set_csum_begin_insert  <= '0';
      set_csum_rsvd_init     <= '0';
      set_txc_addr_0         <= '0';
      set_txc_addr_1         <= '0';
      set_txc_addr_2         <= '0';
      set_txc_addr_3         <= '0';
      set_txc_addr_4_n       <= '0';
      clr_txc_addr_3         <= '0';
      set_txcwr_rd_addr      <= '0';  --  sets the write side, read address to 0x0
      set_txcwr_wr_end       <= '0';  --  writes the end address to the memory in the next available location
      set_txc_en             <= '0';  --  the enable bit to the write side of the memory
      set_txc_we             <= '0';  --  the write enable bit to the write side of the memory
      inc_txd_addr_one       <= '0';
      set_txc_trdy           <= '0';
      init_bram              <= '0';
      compare_addr2          <= '0';
      compare_addr0          <= '0';
      set_txc_trdy2          <= '0';
      clr_txc_trdy2          <= '0';
      enable_compare_addr0_cmplt <= '0';
      inc_txd_addr_one_early <= '0';

      case txc_wr_cs is
        when TXC_ADDR2_WR =>
          set_txc_addr_2         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          txc_wr_ns              <= TXC_ADDR0_WR;
        when TXC_ADDR0_WR =>
          set_txc_addr_0         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          txc_wr_ns              <= WAIT_WR_CMPLT;
        when WAIT_WR_CMPLT =>
          set_txc_addr_0         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          set_txc_trdy2          <= '1';
          txc_wr_ns              <= TXC_WD0;
        when TXC_WD0 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' and
             (wrote_first_packet = '0' or txc_addr_3_dly = '1') then
            set_txc_addr_2         <= '1';  --Set the address to get the TxC Rd Address Pointer
            set_txc_en             <= '1';
            set_axi_flag           <= '1';
            clr_txc_addr_3         <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD1;
          else
            set_txc_addr_2         <= '0';  --Set the address to get the TxC Rd Address Pointer
            set_txc_en             <= '0';
            set_axi_flag           <= '0';
            clr_txc_addr_3         <= '0';
            compare_addr2          <= '0';
            txc_wr_ns              <= TXC_WD0;
          end if;

        when TXC_WD1 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_txc_trdy2          <= '0';
            set_csum_cntrl         <= '1';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD2;--WAIT_ADDR2_COMPARE_CMPLT;
          elsif axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '0' then
          -- need to force txc trdy HIGH since TVALID throttled
            set_txc_trdy2          <= '1';
            set_csum_cntrl         <= '0';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= WAIT_ADDR2_COMPARE_CMPLT;
          else
            set_txc_trdy2          <= '0';
            set_csum_cntrl         <= '0';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD1;
          end if;

        when WAIT_ADDR2_COMPARE_CMPLT =>
        -- now clear txc trdy to only allow a one clock pulse HIGH
          clr_txc_trdy2          <= '1';
          set_txc_addr_2         <= '1';
          set_txc_en             <= '1';
          compare_addr2          <= '1';
          txc_wr_ns              <= TXC_WD1;

        when TXC_WD2 =>
        -- Txc Tready has already been disabled
        --  wait for compare_addr2_cmplt, then
        --  set_txc_trdy2 will force axi_str_txc_tready_int_dly HIGH
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_csum_begin_insert      <= '1';
            set_txc_addr_2         <= '0';
            set_txc_en             <= '0';
            compare_addr2          <= '0';
            set_txc_trdy2          <= '0';
            txc_wr_ns                  <= TXC_WD3;
          else
            if axi_str_txc_tvalid_dly0 = '0'  or
               (txc_mem_full = '1' and axi_str_txc_tvalid_dly0 = '1') then
            --  If full wait for FULL and TVALID
            --  This will allow next elsif to be hit properly
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '1';
              set_txc_en             <= '1';
              compare_addr2          <= '1';
              set_txc_trdy2          <= '0';
              txc_wr_ns              <= TXC_WD2;


            elsif axi_str_txc_tvalid_dly0 = '1' and
              (compare_addr2_cmplt = '1' or compare_addr2_cmplt_dly = '1') then
              --  when full is '0', only need compare_addr2_cmplt to set set_txc_trdy2
              --    which will then allow this state to be exited to TXD_WD3
              --  when full is '1', then will need compare_addr2_cmplt_dly to to set set_txc_trdy2
              --    which will then allow this state to be exited to TXD_WD3
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '0';
              set_txc_en             <= '0';
              compare_addr2          <= '0';
              set_txc_trdy2          <= '1';
              txc_wr_ns                  <= TXC_WD2;
            else
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '1';
              set_txc_en             <= '1';
              compare_addr2          <= '1';
              set_txc_trdy2          <= '0';
              txc_wr_ns                  <= TXC_WD2;
            end if;
          end if;
        when TXC_WD3 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
          --  This is the earliest state to check for TxC FULL from TXC_WD0 state addr_2
          --  Register data, then assert full = 2 clks from rd
          --    Not FULL so write TxC Write Pointer to addr 0x3
            set_csum_rsvd_init         <= '1';
            txc_wr_ns                  <= TXC_WD4;
          else
            set_csum_rsvd_init         <= '0';
            txc_wr_ns                  <= TXC_WD3;
          end if;
        when TXC_WD4 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_txc_addr_0             <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            txc_wr_ns                  <= TXC_WD5;
          else
            set_txc_addr_0             <= '0';  --Set the address to get the TxD Rd Address Pointer
            set_txc_en                 <= '0';
            compare_addr0              <= '0';
            txc_wr_ns                  <= TXC_WD4;
          end if;
        when TXC_WD5 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' and axi_str_txc_tlast_dly0 = '1' then
            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '1';
            txc_wr_ns                  <= WAIT_ADDR0_COMPARE_CMPLT;
          else
            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '0';
            txc_wr_ns                  <= TXC_WD5;
          end if;
        when WAIT_ADDR0_COMPARE_CMPLT =>
          if compare_addr0_cmplt = '1' then
            set_txc_addr_1             <= '1'; -- this is one clock early, so do not set the we enable yet
            set_txc_en                 <= '1';
            set_txc_we                 <= '1';

            set_txc_addr_0             <= '0';
            set_txc_en                 <= '0';
            compare_addr0              <= '0';
            enable_compare_addr0_cmplt <= '0';
            txc_wr_ns                  <= WAIT_TXD_CMPLT;
          else
            set_txc_addr_1             <= '0';
            set_txc_en                 <= '0';
            set_txc_we                 <= '0';

            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '1';
            txc_wr_ns                  <= WAIT_ADDR0_COMPARE_CMPLT;
          end if;



        when WAIT_TXD_CMPLT =>
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1'  and
             axi_str_txd_tlast_dly0 = '1' then
            set_txc_addr_0        <= '0';
            set_txc_addr_1        <= '1';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            if do_csum = '1' then
              inc_txd_addr_one_early <= '1';
            else
              inc_txd_addr_one_early <= '0';
            end if;
            txc_wr_ns             <= WR_TXD_END_PNTR;
          elsif disable_txd_trdy_dly = '1' then
          -- Txd mem is full so get the current read pointer
          --  This can occure after tlast so check it in the following states
            set_txc_addr_0        <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_addr_1        <= '0';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_MEM;
          elsif update_bram_cnt(7) = '1'  then
          --Writing the current TxC write pointer so the read side can monitor it
            set_txc_addr_1        <= '1';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          else
            set_txc_addr_1        <= '0'; --Writing the current TxC write pointer so the read side can monitor it
            set_txc_addr_2        <= '0';
            set_txc_en            <= '0';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          end if;
        when WAIT_TXD_MEM =>
          if disable_txd_trdy_dly = '1' then
            -- Txd mem is full so get the current read pointer
            set_txc_addr_0        <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_addr_1        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_MEM;
          else
            set_txc_addr_0        <= '0';
            set_txc_addr_1        <= '1'; -- this is one clock early, so do not set the we enable yet
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          end if;
        when WR_TXD_END_PNTR =>
          if do_csum = '1' then
            inc_txd_addr_one      <= '1';
            set_txc_addr_4_n      <= '0'; -- Write the TxC End Value to address 0x4 - 0xn
            set_txc_en            <= '0';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_CSUM_END;
          else
            inc_txd_addr_one      <= '1';
            set_txc_addr_4_n      <= '1'; -- Write the TxC End Value to address 0x4 - 0xn
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WR_TXC_PNTR;
          end if;

        when WAIT_CSUM_END =>
          if ptcl_csum_cmplt = '1' then
            inc_txd_addr_one      <= '0'; -- already incremented in WR_TXC_PNTR state
            set_txc_addr_4_n      <= '1'; -- Write the TxC end pointer value to start the tx clint FSM
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WR_TXC_PNTR;
          else
            inc_txd_addr_one      <= '0'; -- already incremented in WR_TXC_PNTR state
            set_txc_addr_4_n      <= '0';
            set_txc_en            <= '0';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_CSUM_END;
          end if;

        when WR_TXC_PNTR =>
          if disable_txc_trdy_dly = '1' then
            set_txc_addr_0        <= '1';
            set_txc_addr_3        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            set_txc_trdy          <= '0';
            txc_wr_ns             <= WR_TXC_PNTR;
          else
            set_txc_addr_0        <= '0'; -- Write the TxC end pointer value to start the tx clint FSM
            set_txc_addr_3        <= '1';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            set_txc_trdy          <= '1';
            txc_wr_ns             <= TXC_WD0;
          end if;

--        when WR_TXC_PNTR =>
--            set_txc_addr_3        <= '1'; -- Write the TxC end pointer value to start the tx clint FSM
--            set_txc_addr_0        <= '0';
--            set_txc_en            <= '1';
--            set_txc_we            <= '1';
--            txc_wr_ns             <= TXC_WD0;

        when others =>
          txc_wr_ns                <= TXC_ADDR2_WR;
      end case;
    end process;

    -----------------------------------------------------------------------------
    -- AXI Stream TX Control State Machine Sequencer
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXC_SEQ : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_wr_cs <= TXC_ADDR2_WR;
        else
          txc_wr_cs <= txc_wr_ns;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    -- Delay the last write to TxC memory of the first packet after reset
    -----------------------------------------------------------------------------
    TX_INIT_INDICATOR_DLYS : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_addr_3_dly2 <= '0';
          txc_addr_3_dly3 <= '0';
        else
          txc_addr_3_dly2 <= txc_addr_3_dly;
          txc_addr_3_dly3 <= txc_addr_3_dly2;
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    -- Use above delay to hold off Tx Client FSM from starting until all
    --    TxD and TxC pointer information has been written to memory
    --
    --    This signal goes through a clock crossing circuit before it is
    --      registered in the Tx Client clock domain and used to start the
    --      Tx Client Read FSM
    -----------------------------------------------------------------------------
    TX_INIT_INDICATOR : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          tx_init_in_prog_int <= '1';
        else
          if txc_addr_3_dly3 = '1' then
            tx_init_in_prog_int <= '0';
          else
            tx_init_in_prog_int <= tx_init_in_prog_int;
          end if;
        end if;
      end if;
    end process;

    tx_init_in_prog <= tx_init_in_prog_int;

    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_1_TXD_WR_PNTR : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_1 = '1' then
          txc_addr_1 <= '1';
        else
          txc_addr_1 <= '0';
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_3_DELAY : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' or clr_txc_addr_3 = '1' then
          txc_addr_3_dly  <= '0';
        elsif set_txc_addr_3 = '1' then
          txc_addr_3_dly <= '1';
        else
          txc_addr_3_dly <= txc_addr_3_dly;
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    --  Generate address that will hold the End Address
    -----------------------------------------------------------------------------
    TXC_WR_ADDR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_mem_wr_addr      <= txc_min_wr_addr;
          txc_mem_wr_addr_last <= txc_wr_addr3;
          txc_mem_wr_addr_0    <= txc_wr_addr5;
          txc_mem_wr_addr_1    <= txc_wr_addr6;
        else
          if set_txc_addr_3 = '1' then
            --  increment the address for the next packet
            --  use the delayed signal to increment after the current address
            --  can be written
            if txc_mem_wr_addr = txc_max_wr_addr then
              --  if the max address is reached, loop to address 0x4
              txc_mem_wr_addr      <= txc_mem_wr_addr_0;
              txc_mem_wr_addr_last <= txc_wr_addr3;
              txc_mem_wr_addr_0    <= txc_mem_wr_addr_1;  --plus1
              txc_mem_wr_addr_1    <= txc_wr_addr6;       --plus2
            else
              --  otherwise just increment it
              txc_mem_wr_addr      <= txc_mem_wr_addr_0;
              txc_mem_wr_addr_last <= txc_mem_wr_addr;
              txc_mem_wr_addr_0    <= txc_mem_wr_addr_1;
              txc_mem_wr_addr_1    <= std_logic_vector(unsigned(txc_mem_wr_addr_1) + 1);
            end if;
          else -- Hold the current address until something changes
            txc_mem_wr_addr      <= txc_mem_wr_addr;
            txc_mem_wr_addr_last <= txc_mem_wr_addr_last;
            txc_mem_wr_addr_0    <= txc_mem_wr_addr_0;
            txc_mem_wr_addr_1    <= txc_mem_wr_addr_1;
          end if;
        end if;
      end if;
    end process;




    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_0_DELAY : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        txc_addr_0_dly1 <= set_txc_addr_0;
        txc_addr_0_dly2 <= txc_addr_0_dly1;
      end if;

    end process;


    -----------------------------------------------------------------------------
    --  Generate address that will hold the End Address
    -----------------------------------------------------------------------------
    MEM_TXC_WR_ADDR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then

        if set_txc_addr_4_n = '1' and set_txc_we = '1' then
          -- Provide the address for the End of packet address
          Axi_Str_TxC_2_Mem_Addr_int <= txc_mem_wr_addr;
        elsif set_txc_addr_3 = '1' and set_txc_we = '1' then
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr3; --set txc wr pointer
        elsif txc_addr_2 = '1' and  (txc_we = '0' or init_bram = '1') then
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr2; --get txc rd pointer
        elsif set_txc_addr_0 = '1' and (set_txc_we = '0' or init_bram = '1') then
          --  Monitor the read pointer for a full
          --  condition in the TxD Memory
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr0;
        elsif set_txc_addr_1 = '1' then
          --  Set the TxD write pointer to
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr1;
        else
          Axi_Str_TxC_2_Mem_Addr_int <= (others => '0');
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_Addr <= Axi_Str_TxC_2_Mem_Addr_int;
    txc_mem_wr_addr_plus1  <= txc_mem_wr_addr_0;
    txc_mem_wr_addr_plus2  <= txc_mem_wr_addr_1;

    -----------------------------------------------------------------------------
    --  This process remaps the strobe signal to the byte address offset minus
    --  one byte.
    -----------------------------------------------------------------------------
    END_ADDRESS_BYTE_OFFSET : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txD = '1' then
          end_addr_byte_offset <= (others => '0');
        elsif axi_str_txd_tlast_dly0 = '1' and axi_str_txd_tvalid_dly0 = '1' and
              axi_str_txd_tready_int_dly = '1' then
          case axi_str_txd_tstrb_dly0 is
            when "1111" => end_addr_byte_offset <= "11";
            when "0111" => end_addr_byte_offset <= "10";
            when "0011" => end_addr_byte_offset <= "01";
            when others => end_addr_byte_offset <= "00";
          end case;
        else
          end_addr_byte_offset <= end_addr_byte_offset;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_WR_ADDR_VALUE : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' or init_bram = '1' then
          Axi_Str_TxC_2_Mem_Din_int <= (others => '0');

        elsif set_txc_addr_4_n = '1' and do_csum = '0' then
        --write the ending address of the packet to memory minus one byte
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd_2 & axi_str_txd_2_mem_addr_int & end_addr_byte_offset;
        elsif set_txc_addr_4_n = '1' and do_csum = '1' then
        -- Increment already happened so use current value
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd_2 & axi_str_txd_2_mem_addr_int_mins1 & end_addr_byte_offset;
        elsif set_txc_addr_3 = '1' then
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txc & txc_mem_wr_addr;
        else
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd & axi_str_txd_2_mem_addr_int_plus1;
        end if;
      end if;
    end process;



    Axi_Str_TxC_2_Mem_Din <= Axi_Str_TxC_2_Mem_Din_int;

  --  Axi_Str_TxC_2_Mem_En  <= '1';
    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if (set_txc_en = '1' and set_txc_addr_2 = '0') or
           addr_2_en = '1' or init_bram = '1' then
          Axi_Str_TxC_2_Mem_En <= '1';
        else
          Axi_Str_TxC_2_Mem_En <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_WR_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_we = '1' then
          Axi_Str_TxC_2_Mem_We_int(0) <= '1';
        else
          Axi_Str_TxC_2_Mem_We_int(0) <= '0';
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_We <= Axi_Str_TxC_2_Mem_We_int;


    -----------------------------------------------------------------------------
    --  Delay set_txc_addr_2 to align with data
    -----------------------------------------------------------------------------
    TXC_ADDR2_DLY : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_2 = '1' then
          txc_addr_2  <= set_txc_addr_2;
        else
          txc_addr_2  <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay set_txc_we to align with address
    -----------------------------------------------------------------------------
    TXC_WE_DLY : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_we = '1' then
          txc_we  <= set_txc_we;
        else
          txc_we  <= '0';
        end if;
        txc_we_dly1 <= txc_we;
        txc_we_dly2 <= txc_we_dly1;

      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay set_txc_we to align with address
    -----------------------------------------------------------------------------
    ADDR2_MEM_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_2 = '1' and  set_txc_en = '1' then
          addr_2_en  <= set_txc_en;
        else
          addr_2_en  <= '0';
        end if;
        addr_2_en_dly1 <= addr_2_en;
        addr_2_en_dly2 <= addr_2_en_dly1;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Get the read pointer to check for FULL
    --  With ASYNC BRAM clock cannot read/write same address in memory at same
    --  time unless timing is met, so read until data matches
    -----------------------------------------------------------------------------
    MEM_TXC_RD_ADDR_PNTR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_rd_addr2_pntr_1 <= (others => '0');
          txc_rd_addr2_pntr   <= txc_min_wr_addr;
          compare_addr2_cmplt <= '0';
          compare_addr2_cmplt_dly <= '0';
        else

          if set_txc_addr_2 = '1' and addr_2_en_dly2 = '1' and txc_we_dly2 = '0' then
            txc_rd_addr2_pntr_1 <= Axi_Str_TxC_2_Mem_Dout(c_TxC_addrb_width -1 downto 0);

            if Axi_Str_TxC_2_Mem_Dout(c_TxC_addrb_width -1 downto 0) = txc_rd_addr2_pntr_1  and
               compare_addr2_cmplt = '0' then
              txc_rd_addr2_pntr   <= txc_rd_addr2_pntr_1;
              compare_addr2_cmplt <= '1';
            else
              txc_rd_addr2_pntr   <= txc_rd_addr2_pntr;
              compare_addr2_cmplt <= '0';
            end if;

          else
            txc_rd_addr2_pntr_1 <= txc_rd_addr2_pntr_1;
            txc_rd_addr2_pntr   <= txc_rd_addr2_pntr;
            compare_addr2_cmplt <= '0';
          end if;
          compare_addr2_cmplt_dly <= compare_addr2_cmplt;

        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Full flag indicator
    --    Does not begin comparison until 1st packet is written to memory
    -----------------------------------------------------------------------------
    TXC_FULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txc = '1' then
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
        elsif txc_mem_full = '1' and
           compare_addr2_cmplt = '1' and compare_addr2_cmplt_dly = '0' then
           --increments after it goes full, so use txc_mem_wr_addr for compare
          if txc_mem_wr_addr /= txc_rd_addr2_pntr then
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
          else
            txc_mem_full     <= txc_mem_full;
            txc_mem_not_full <= txc_mem_not_full;
          end if;
        elsif set_txc_addr_3 = '1' and set_txc_we = '1' then
          if txc_mem_wr_addr_plus1 = txc_rd_addr2_pntr then
            txc_mem_full     <= '1';
            txc_mem_not_full <= '0';
          else
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
          end if;
        else
          txc_mem_full     <= txc_mem_full;
          txc_mem_not_full <= txc_mem_not_full;
        end if;
      end if;
    end process;

    TXC_AFULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if txc_mem_wr_addr_plus2 = txc_rd_addr2_pntr then
          txc_mem_afull     <= '1';
        else
          txc_mem_afull     <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Throttle AXI Stream TxC
    --    Do not assert unless TxD is not in progress and the memory can
    --    accept data
    -----------------------------------------------------------------------------
    TXC_READY : process(AXI_STR_TXD_ACLK)
    begin



      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txc = '1' or clr_txc_trdy = '1' or clr_txc_trdy2 = '1' or
             set_txd_rdy = '1' or (txd_rdy = '1' and clr_txd_rdy = '0') or disable_txc_trdy = '1' or
             (AXI_STR_TXC_TLAST = '1' and AXI_STR_TXC_TVALID = '1' and axi_str_txc_tready_int = '1') or
             (compare_addr2 = '1' and axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1') then --do not need compare_addr0 because will clr at TLAST
          axi_str_txc_tready_int <= '0';
        else

          if txc_addr_3_dly = '1' then
            if (txc_mem_wr_addr = txc_rd_addr2_pntr and txc_mem_full = '1') then
              axi_str_txc_tready_int <= '0';
            elsif txc_mem_wr_addr = txc_rd_addr2_pntr and
                Axi_Str_TxC_2_Mem_We_int(0) = '1' then
              axi_str_txc_tready_int <= '0';
            else
              axi_str_txc_tready_int <= axi_str_txc_tready_int;
            end if;
          elsif set_txc_trdy = '1' then
            axi_str_txc_tready_int <= '1';
          elsif set_txc_trdy2 = '1' then
          --  need to force it high after address compare and after reset
            axi_str_txc_tready_int <= '1';
          else
            axi_str_txc_tready_int <= axi_str_txc_tready_int;
          end if;
        end if;
        axi_str_txc_tready_int_dly <= axi_str_txc_tready_int;
      end if;
    end process;

    AXI_STR_TXC_TREADY <= axi_str_txc_tready_int;

    -----------------------------------------------------------------------------
    --  Register and hold the axi_flag information and CSUM Control information
    --    axi_flag
    --      0x5 = Status control
    --      0xA = Normal control
    --      0xF = Null Control
    --    CSUM
    --      00 = No CSUM will be performed
    --      01 = Partial Checksum will be performed
    --      10 = Full checksum offloading will be performed
    -----------------------------------------------------------------------------
    CNTRL_WD0 : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          axi_flag   <= (others => '0');
        elsif set_axi_flag = '1' then
          axi_flag   <= axi_str_txc_tdata_dly0(31 downto 28);
        else
          axi_flag   <= axi_flag;
        end if;
      end if;
    end process;

    CNTRL_WD1 : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          csum_cntrl <= (others => '0');
        elsif set_csum_cntrl = '1' then
          csum_cntrl <= axi_str_txc_tdata_dly0 (1 downto  0);
        else
          csum_cntrl <= csum_cntrl;
        end if;
      end if;
    end process;

      ---------------------------------------------------------------------------
      --  Delay signal to load csum value in csum calculation
      ---------------------------------------------------------------------------
      CHECK_FULL_SIG : process(AXI_STR_TXC_ACLK)
      begin

        if rising_edge(AXI_STR_TXC_ACLK) then
          check_full <= set_txc_addr_4_n;
        end if;
      end process;


    -----------------------------------------------------------------------------
    --  This generate is used to reduce a small amount of logic when the CSUM
    --    functionality is not included in the build
    -----------------------------------------------------------------------------
    GEN_CSUM_SUPPORT : if C_TXCSUM = 2 generate
    begin

      ---------------------------------------------------------------------------
      --  Store the starting address of the frame which is used to calculate
      --  the address where the IPv4 Header CSUM and the TCP/UDP header CSUM
      --  will be written in BRAM memory
      ---------------------------------------------------------------------------
      CSUM_START_ADDR : process(AXI_STR_TXC_ACLK)
      begin

        if rising_edge(AXI_STR_TXC_ACLK) then
          if reset2axi_str_txc = '1' or clr_csums = '1' then
            csum_strt_addr <= (others => '0');
          else
            if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' and
               axi_str_txc_tlast_dly0 = '1' then
               csum_strt_addr <= axi_str_txd_2_mem_addr_int;
            else
               csum_strt_addr <= csum_strt_addr;
            end if;
          end if;
        end if;
      end process;

      ---------------------------------------------------------------------
      --  Use the FLAG field in the TxC AXI Stream to enable the CSUM on
      --  a frame by frame basis if needed.  This will stay set until the
      --  flag on the following frame unsets it, or if all of the criteria
      --  for the Full CSUM is not met and the calculation is aborted.
      --
      --  This signal is used in conjunction with ptcl_csum_cmplt to allow
      --  the CSUM calculation to be written to the memory when all of the
      --  CSUM criteria has been met.
      ---------------------------------------------------------------------
      CSUM_ENABLE : process(AXI_STR_TXC_ACLK)
      begin

        if rising_edge(AXI_STR_TXC_ACLK) then
--          if reset2axi_str_txc = '1' or abort_csum = '1' then
          --  if any of the requirements to perform a full csum are not met,
          --  the FSM will exit early, so clear this signal
          if reset2axi_str_txc = '1' then
          --  Originally used abort_csum to clear when FULL_CSUM_FSM_TYPE returned to idle before end of packet
          --  Changed FSM to wait until after end of packet and return to idle with other FSMs
            do_csum <= '0';
          else
            if axi_str_txc_tready_int_dly = '1' and
               axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tlast_dly0 = '1' then
              case axi_flag is
                when "1010" =>
                  case csum_cntrl is
                    when "10"   => do_csum <= '1';
                    when others => do_csum <= '0';
                  end case;
                when others =>
                  do_csum <= '0';
              end case;
            else
              do_csum <= do_csum;
            end if;
          end if;
        end if;
      end process;


      csum_calc_en  <= axi_str_txd_tvalid_dly0 and axi_str_txd_tready_int_dly;


      I_TX_FCSUM_HDR_CALC : tx_csum_full_calc_if
      generic map(
        C_IPV4_HEADER_CSUM => 1
      )
      port map (
        clk               => AXI_STR_TXD_ACLK,
        reset             => reset2axi_str_txd,
        clr_csums         => clr_csums,
        txd_tlast         => axi_str_txd_tlast_dly0,
        csum_calc_en      => csum_calc_en,

        tcp_ptcl          => tcp_ptcl,
        udp_ptcl          => udp_ptcl,
        do_ipv4hdr        => do_ipv4hdr,
        not_tcp_udp       => not_tcp_udp,
        do_full_csum      => do_full_csum,

        do_csum           => do_csum,
        csum_en_b32       => en_ipv4_hdr_b32,
        csum_en_b10       => en_ipv4_hdr_b10,
        zeroes_en         => zeroes_en,

        data_last         => last_ipv4_hdr_cnt,
        inc_txd_addr_one  => inc_txd_addr_one,
        inc_txd_addr_one_early => inc_txd_addr_one_early,

        csum_din          => csum_din,
        csum_dout         => hdr_csum_dout,
        csum_we           => hdr_csum_we,       -- not used  (comb)
        csum_cmplt        => hdr_csum_cmplt

      );

      I_TX_FCSUM_DATA_CALC : tx_csum_full_calc_if
      generic map(
        C_IPV4_HEADER_CSUM => 0
      )
      port map (
        clk               => AXI_STR_TXD_ACLK,
        reset             => reset2axi_str_txd,
        clr_csums         => clr_csums,
        txd_tlast         => axi_str_txd_tlast_dly0,
        csum_calc_en      => csum_calc_en,

        tcp_ptcl          => tcp_ptcl,
        udp_ptcl          => udp_ptcl,
        do_ipv4hdr        => do_ipv4hdr,
        not_tcp_udp       => not_tcp_udp,
        do_full_csum      => do_full_csum,

        do_csum           => do_csum,
        csum_en_b32       => fsm_csum_en_b32,
        csum_en_b10       => fsm_csum_en_b10,
        zeroes_en         => zeroes_en,

        data_last         => add_psdo_wd,
        inc_txd_addr_one  => inc_txd_addr_one,
        inc_txd_addr_one_early => inc_txd_addr_one_early,

        csum_din          => csum_din,
        csum_dout         => ptcl_csum_dout,
        csum_we           => ptcl_csum_we,      -- not used (comb)
        csum_cmplt        => ptcl_csum_cmplt    -- this always pulses for one clock
      );                                        -- whether or not the CSUM was calculated or not
                                                -- It is used to allow the Txc FSM to sequence back to
                                                -- to its starting state for the next packet and also
                                                -- in conjunction with do_csum to write the memory with
                                                -- the csum calculation when the Full CSUM is calculated


      I_TX_FULL_CSUM_FSM : tx_csum_full_fsm
      generic map(
        C_S_AXI_DATA_WIDTH  => C_S_AXI_DATA_WIDTH,
        c_TxD_addrb_width   => c_TxD_addrb_width
      )
      port map(

        AXI_STR_TXD_ACLK  => AXI_STR_TXD_ACLK,
        reset2axi_str_txd => reset2axi_str_txd,

        txd_strbs         => axi_str_txd_tstrb_dly0,
        do_csum           => do_csum,           -- : in  std_logic;  --  axi_flag must = 0xA for this to be enabled
        abort_csum        => abort_csum,        -- : out std_logic;  -: out std_logic;  -
        txd_tlast         => axi_str_txd_tlast_dly0, -- : in  std_logic;
        csum_calc_en      => csum_calc_en,      -- : in  std_logic;  --  axi_str_txd_tvalid_dly0 and axi_str_txd_tready_int_dly;
        clr_csums         => clr_csums,         -- : out std_logic;  --  Clear CSUM flags and calculations
        tcp_ptcl          => tcp_ptcl,          -- : out std_logic;  --  TCP Protocol Indicator
        udp_ptcl          => udp_ptcl,          -- : out std_logic;  --  UDP Protocol Indicator
        en_ipv4_hdr_b32   => en_ipv4_hdr_b32,   -- : out std_logic_vector( 1 downto 0);  --  bytes 3 and 2 of din
        en_ipv4_hdr_b10   => en_ipv4_hdr_b10,   -- : out std_logic_vector( 1 downto 0);  --  bytes 1 and 0 of din
        last_ipv4_hdr_cnt => last_ipv4_hdr_cnt, -- : out std_logic;                      --  last data for IPv4 Header Calculation
        fsm_csum_en_b32   => fsm_csum_en_b32,   -- : out std_logic_vector( 1 downto 0);  --  bytes 3 and 2 of din
        fsm_csum_en_b10   => fsm_csum_en_b10,   -- : out std_logic_vector( 1 downto 0);  --  bytes 1 and 0 of din
        add_psdo_wd       => add_psdo_wd,       -- : out std_logic;                      --  last data for TCP/UDP Calculation
        ptcl_csum_cmplt   => ptcl_csum_cmplt,   -- : in  std_logic;                      --  indicates the TCP/UDP csum calculation is complete or used to finish a non-csum frame
        zeroes_en         => zeroes_en,         -- : out std_logic_vector( 1 downto 0);  --  stalls the CSUM calculations for one clock so Zeroes do not need muxed in
        din               => axi_str_txd_tdata_dly0, -- : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1  downto 0) -- AXI Stream Tx Data
        csum_din          => csum_din,          -- : out std_logic_vector(C_S_AXI_DATA_WIDTH-1  downto 0) -- mux out
        do_ipv4hdr        => do_ipv4hdr,      -- out std_logic
        not_tcp_udp       => not_tcp_udp,    --: out std_logic;      --  only do the ipv4 header csum - no TCP/UDP protocol

        do_full_csum      => do_full_csum,    -- out std_logic
        hdr_csum_cmplt    => hdr_csum_cmplt,
        wr_hdr_csum       => wr_hdr_csum,       -- : out std_logic
        wr_ptcl_csum      => wr_ptcl_csum,      -- : out std_logic

        csum_strt_addr    => csum_strt_addr,    -- : in  std_logic_vector(c_TxD_addrb_width-1   downto 0);starting address of the packet
        csum_ipv4_hdr_addr=> csum_ipv4_hdr_addr,-- : out std_logic_vector(c_TxD_addrb_width-1   downto 0);
        csum_ipv4_hdr_we  => csum_ipv4_hdr_we,  -- : out std_logic_vector( 3 downto 0);
        csum_ptcl_addr    => csum_ptcl_addr,    -- : out std_logic_vector(c_TxD_addrb_width-1   downto 0);
        csum_ptcl_we      => csum_ptcl_we       -- : out std_logic_vector( 3 downto 0)
      );

    end generate GEN_CSUM_SUPPORT;


    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Data Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXD_CONTROL : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_tvalid_dly0 <= '0';
          axi_str_txd_tlast_dly0  <= '0';
          clr_txd_trdy            <= '0';
        else
          axi_str_txd_tvalid_dly0 <= AXI_STR_TXD_TVALID;
          axi_str_txd_tlast_dly0  <= AXI_STR_TXD_TLAST;
          if axi_str_txd_tvalid = '1' and axi_str_txd_tlast = '1' and axi_str_txd_tready_int = '1' then
            clr_txd_trdy <= '1';
          else
            clr_txd_trdy <= '0';
          end if;
        end if;
      end if;
    end process;

    AXI_STR_TXD_TREADY <= axi_str_txd_tready_int;  --fix me  need to look at all txd control and TXC tlast

    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Data Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXD_IN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_tstrb_dly0  <= AXI_STR_TXD_TSTRB;
        axi_str_txd_tdata_dly0  <= AXI_STR_TXD_TDATA;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Delay the data one more clock for BRAM
    -----------------------------------------------------------------------------
    REG_TXD_DLY0 : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
          if wr_hdr_csum = '1' then
          -- Mux in the CSUM result
            --  The WE will only allow a 16 bit write to memory
            axi_str_txd_tdata_dly1 <= hdr_csum_dout & hdr_csum_dout;
          elsif ptcl_csum_cmplt = '1' and do_full_csum = '1'  then
          -- Write the memory with the csum calculation
          -- Mux in the CSUM result
            --  The WE will only allow a 16 bit write to memory
            axi_str_txd_tdata_dly1 <= ptcl_csum_dout & ptcl_csum_dout;
          elsif axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
            axi_str_txd_tdata_dly1  <= axi_str_txd_tdata_dly0;
          else
            axi_str_txd_tdata_dly1  <= axi_str_txd_tdata_dly1;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  AXI Stream TX Data State Machine - combinational/combinatorial
    --    Used to provide the control to write the data to the BRAM
    --    This state machine will throttle the Transmit AXI Stream Control state
    --      machine until after the data information has been received.
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXD_CMB : process (txd_wr_cs,axi_str_txd_tvalid_dly0,
      axi_str_txd_tlast_dly0,
      axi_str_txd_tstrb_dly0,wrote_first_packet,axi_str_txd_tready_int_dly,
      txd_rd_pntr,txd_mem_full,txd_min_wr_addr,
      txd_rd_pntr_hold,do_csum,txd_rdy,ptcl_csum_cmplt,txd_mem_afull,txd_rd_pntr_hold_plus3,
      compare_addr0_cmplt,do_ipv4hdr,do_full_csum,
      axi_str_txd_2_mem_addr_int,txd_max_wr_addr,
      check_full,txd_max_wr_addr_minus4)
    begin

      inc_txd_wr_addr     <= '0';
      set_txd_we          <= "0000";
      set_txd_en          <= '0';
      set_first_packet    <= '0';
      set_txd_rdy         <= '0';
      clr_txd_rdy         <= '0';
      clr_full_pntr       <= '0';
      disable_txd_trdy    <= '0';
      disable_txc_trdy    <= '0';
      halt_pntr_update    <= '0';
      set_txd_mem_full    <= '0';
      clr_txd_mem_full    <= '0';
      set_txd_mem_afull   <= '0';
      update_rd_pntrs     <= '0';

      case txd_wr_cs is
        when IDLE =>
          if compare_addr0_cmplt = '1' then
          --  Requirement is that the TXD and TXC interfaces use the same clock
          --    so it is OK to used the TXC signals in the TXD state machine
            set_txd_rdy <= '1';
            txd_wr_ns   <= TXD_PRM;
          else
            set_txd_rdy <= '0';
            txd_wr_ns   <= IDLE;
          end if;
        when TXD_PRM =>
--      Made change to ensure TxD Memory is never full here.
--      The memory can always accept data at the start of a transfer
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
          --  delay incrementing pointer until next data
          --    Ethernet has to send 14bytes as a bare minimum, so it is
          --    guaranteed to get through this state with all of the strobes set
          --    and TLAST = '0'
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            disable_txd_trdy    <= '0';
            txd_wr_ns           <= TXD_WRT;
          else
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            disable_txd_trdy    <= '0';
            txd_wr_ns           <= TXD_PRM;
          end if;
        when  TXD_WRT =>
          if txd_mem_full = '1' and axi_str_txd_tready_int_dly = '0' then
          --memory is full when axi_str_txd_tready_int_dly = '0'
            inc_txd_wr_addr     <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_first_packet    <= '0';
            clr_txd_rdy         <= '0';
            disable_txd_trdy    <= '1';
            txd_wr_ns           <= MEM_FULL;
          elsif axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
            inc_txd_wr_addr     <= '1';
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            if axi_str_txd_tlast_dly0 = '1' then
              if do_csum = '1' then
              --  do not care if memory is full because we are over-writing
              --  a location
                set_first_packet    <= '0';
                clr_txd_rdy         <= '1';
                disable_txc_trdy    <= '1';
                disable_txd_trdy    <= '0';
                txd_wr_ns           <= WAIT_CSUM;
              else-- txd_mem_full = '1' or txd_mem_afull = '1'
              --  received TLAST but fifo is full so wait until it can
              --  accept more data before going idle

                if wrote_first_packet = '0' then
                  set_first_packet <= '1';
                else
                  set_first_packet <= '0';
                end if;

                clr_txd_rdy         <= '1';
                disable_txc_trdy    <= '1';
                disable_txd_trdy    <= '0';
                txd_wr_ns           <= WAIT_WR1;
              end if;
            else
            --  received data (normal receive), so continue receiving data
              set_first_packet    <= '0';
              clr_txd_rdy         <= '0';
              disable_txd_trdy    <= '0';
              txd_wr_ns           <= TXD_WRT;
            end if;
          else
            inc_txd_wr_addr     <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_first_packet    <= '0';
            clr_txd_rdy         <= '0';
            disable_txd_trdy    <= '0';
            txd_wr_ns           <= TXD_WRT;
          end if;
       when MEM_FULL =>
          --  stay here until the read pointer updates by 4 words or more.  The read side operates on bytes,
          --  the write side operates on words.
          --    The read pointer updates every 512 bytes (128 words) and at the end of a packet.
          --      The samallest packet the can be sent is 15bytes, but since the BRAM is 32 bit aligned,
          --      the read side will usually update the read pointer by a minimum of 16 bytes (4 words).  However,
          --      it can update by by less than 16 bytes (4 words).  This can occure if a packet started at read
          --      address 0x1A4 (write address 0x69), and the packet is 516 bytes in length (129 words).  Here the read pointer
          --      will update at 0x3A4 (write address 0xE9 - 128 words) then again at the end of the packet at 0x3A8
          --      (write address 0xEA).
          --        If this occures the below logic will detect it and update the read pointer, but stay in this
          --        state until the next update occurs.  The next update is guaranteed to be greater than 4 words,
          --        which will allow the full pointers to be cleared for the next packet.
          inc_txd_wr_addr     <= '0';
          set_txd_we          <= "0000";
          set_txd_en          <= '0';
          set_first_packet    <= '0';
          clr_txd_rdy         <= '0';
          if txd_rd_pntr = txd_rd_pntr_hold then
          --  stay here until an update occurs
            update_rd_pntrs  <= '0';
            disable_txd_trdy <= '1';
            clr_full_pntr    <= '0';
            txd_wr_ns        <= MEM_FULL;
          else
          --  The read pointer was updated to determine if it was updated by 4 words or more
          --    If not, update the hold pointers, but stay in this state
            if txd_rd_pntr_hold <= txd_max_wr_addr_minus4 then
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x0 - 0x1FB
              if txd_rd_pntr > txd_rd_pntr_hold_plus3 then
              -- an update of 4 words or greater occured so exit this state
                update_rd_pntrs  <= '0';
                disable_txd_trdy <= '0';
                clr_full_pntr    <= '1';
                txd_wr_ns        <= TXD_WRT;
              else
              --  the update was less than 4 words
              --    (txd_rd_pntr <= txd_rd_pntr_hold_plus3)
                if txd_rd_pntr < txd_rd_pntr_hold then
                --  the read pointer wrapped, so exit because the update was > 4 words
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              end if;
            else
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x1FC- 0x1FF
              if txd_rd_pntr_hold_plus3 = txd_max_wr_addr then
              --  txd_rd_pntr = 0x1FC for 2048 byte memory, so txd_rd_pntr_hold_plus3 = max memory size
                if (txd_rd_pntr <= txd_rd_pntr_hold) then
                --  the update was >= 4 words so exit
                --    for a 2048 memory, txd_rd_pntr_hold = 0x1FC
                --      if txd_rd_pntr is between 0x0 and 0x1FB then an update of 4 or more words occurred
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              else
              --  txd_rd_pntr = 0x1FD, 0x1FE, or 0x1FF for 2048 byte memory,
              --  so the minimum txd_rd_pntr_hold_plus3 can be is 0, 1, or 2
                if (txd_rd_pntr > txd_rd_pntr_hold_plus3) and (txd_rd_pntr < txd_rd_pntr_hold) then
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr has to be tween 0x1 and 0x1FC to exit this state
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr has to be tween 0x2 and 0x1FD to exit this state
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr has to be tween 0x3 and 0x1FE to exit this state
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  txd_rd_pntr did not update by 4 or more words, so update hold poointers and stay in this state
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited BUT
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr was only updated 1-3 words to 0x1FE, 0x1FF, or 0x0, so stay here
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr was only updated 1-3 words to 0x1FF, 0x0, or 0x1, so stay here
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr was only updated 1-3 words to 0x0, 0x1, or 0x2, so stay here
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              end if;
            end if;
          end if;

        when CLR_FULL =>
          --  stay here until the read pointer updates by 4 words or more.  The read side operates on bytes,
          --  the write side operates on words.
          --    The read pointer updates every 512 bytes (128 words) and at the end of a packet.
          --      The samallest packet the can be sent is 15bytes, but since the BRAM is 32 bit aligned,
          --      the read side will usually update the read pointer by a minimum of 16 bytes (4 words).  However,
          --      it can update by by less than 16 bytes (4 words).  This can occure if a packet started at read
          --      address 0x1A4 (write address 0x69), and the packet is 516 bytes in length (129 words).  Here the read pointer
          --      will update at 0x3A4 (write address 0xE9 - 128 words) then again at the end of the packet at 0x3A8
          --      (write address 0xEA).
          --        If this occures the below logic will detect it and update the read pointer, but stay in this
          --        state until the next update occurs.  The next update is guaranteed to be greater than 4 words,
          --        which will allow the full pointers to be cleared for the next packet.
          inc_txd_wr_addr     <= '0';
          set_txd_we          <= "0000";
          set_txd_en          <= '0';
          set_first_packet    <= '0';
          clr_txd_rdy         <= '0';
          if txd_rd_pntr = txd_rd_pntr_hold then
          --  stay here until an update occurs
            update_rd_pntrs  <= '0';
            halt_pntr_update <= '1';
            disable_txc_trdy <= '1';
            disable_txd_trdy <= '1';
            clr_full_pntr    <= '0';
            txd_wr_ns        <= CLR_FULL;
          else
          --  The read pointer was updated to determine if it was updated by 4 words or more
          --    If not, update the hold pointers, but stay in this state
            if txd_rd_pntr_hold <= txd_max_wr_addr_minus4 then
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x0 - 0x1FB
              if txd_rd_pntr > txd_rd_pntr_hold_plus3 then
              -- an update of 4 words or greater occured so exit this state
                if wrote_first_packet = '0' then
                  set_first_packet <= '1';
                else
                  set_first_packet <= '0';
                end if;
                update_rd_pntrs  <= '0';
                halt_pntr_update <= '0';
                disable_txd_trdy <= '0';
                clr_full_pntr    <= '1';
                clr_txd_rdy      <= '0';
                txd_wr_ns        <= WAIT_COMPARE_CMPLT;
              else
              --  the update was less than 4 words
              --    (txd_rd_pntr <= txd_rd_pntr_hold_plus3)
                if txd_rd_pntr < txd_rd_pntr_hold then
                --  the read pointer wrapped, so exit because the update was > 4 words
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  halt_pntr_update <= '1';
                  disable_txc_trdy <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= CLR_FULL;
                end if;
              end if;
            else
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x1FC- 0x1FF
              if txd_rd_pntr_hold_plus3 = txd_max_wr_addr then
              --  txd_rd_pntr = 0x1FC for 2048 byte memory, so txd_rd_pntr_hold_plus3 = max memory size
                if (txd_rd_pntr <= txd_rd_pntr_hold) then
                --  the update was >= 4 words so exit
                --    for a 2048 memory, txd_rd_pntr_hold = 0x1FC
                --      if txd_rd_pntr is between 0x0 and 0x1FB then an update of 4 or more words occurred
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  halt_pntr_update <= '1';
                  disable_txc_trdy <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= CLR_FULL;
                end if;
              else
              --  txd_rd_pntr = 0x1FD, 0x1FE, or 0x1FF for 2048 byte memory,
              --  so the minimum txd_rd_pntr_hold_plus3 can be is 0, 1, or 2
                if (txd_rd_pntr > txd_rd_pntr_hold_plus3) and (txd_rd_pntr < txd_rd_pntr_hold) then
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr has to be tween 0x1 and 0x1FC to exit this state
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr has to be tween 0x2 and 0x1FD to exit this state
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr has to be tween 0x3 and 0x1FE to exit this state
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  txd_rd_pntr did not update by 4 or more words, so update hold poointers and stay in this state
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited BUT
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr was only updated 1-3 words to 0x1FE, 0x1FF, or 0x0, so stay here
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr was only updated 1-3 words to 0x1FF, 0x0, or 0x1, so stay here
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr was only updated 1-3 words to 0x0, 0x1, or 0x2, so stay here
                  update_rd_pntrs  <= '1';
                  halt_pntr_update <= '1';
                  disable_txc_trdy <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= CLR_FULL;
                end if;
              end if;
            end if;
          end if;
        when WAIT_CSUM =>
          if txd_mem_full = '1' then -- hold until complete with CSUM
            set_txd_mem_full <= '1';
          else
            set_txd_mem_full <= '0';
          end if;

          if txd_mem_afull = '1' then -- hold until complete with CSUM
            set_txd_mem_afull <= '1';
          else
            set_txd_mem_afull <= '0';
          end if;

          if ptcl_csum_cmplt = '1' then --one clock cycle pulse
            if txd_mem_full = '1' or txd_mem_afull = '1' then
              set_first_packet  <= '0';
              disable_txc_trdy  <= '1';
              disable_txd_trdy  <= '1';
              clr_txd_mem_full  <= '0';
              txd_wr_ns         <= CLR_FULL;
            else
              if wrote_first_packet = '0' then
                set_first_packet <= '1';
              else
                set_first_packet <= '0';
              end if;
              set_first_packet  <= '0';
              disable_txc_trdy  <= '0';
              disable_txd_trdy  <= '0';
              clr_txd_mem_full  <= '0';
              txd_wr_ns         <= IDLE;
            end if;
          else
            clr_txd_rdy       <= '0';
            disable_txc_trdy  <= '1';
            clr_txd_mem_full  <= '0';
            txd_wr_ns         <= WAIT_CSUM;
          end if;

        when WAIT_WR1 =>
          disable_txc_trdy  <= '1';
          disable_txd_trdy  <= '0';

          if check_full = '1' then
            txd_wr_ns         <= WAIT_WR2;
          else
            txd_wr_ns         <= WAIT_WR1;
          end if;
        when WAIT_WR2 =>
          if txd_mem_full = '1' or txd_mem_afull = '1' then
            disable_txc_trdy  <= '1';
            disable_txd_trdy  <= '1';
            txd_wr_ns         <= CLR_FULL;
          else
            if wrote_first_packet = '0' then
              set_first_packet <= '1';
            else
              set_first_packet <= '0';
            end if;

            disable_txc_trdy  <= '0';
            disable_txd_trdy  <= '0';
            txd_wr_ns         <= IDLE;
          end if;
        when WAIT_COMPARE_CMPLT =>
          txd_wr_ns        <= IDLE;
        when others =>
          txd_wr_ns <= IDLE;
      end case;
    end process;

    -----------------------------------------------------------------------------
    -- AXI Stream TX Control State Machine Sequencer
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXD_SEQ : process (AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_wr_cs <= IDLE;
        else
          txd_wr_cs <= txd_wr_ns;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    -- Indicator when performing a write to TxD Memory
    --  clear on axi_str_txd_tlast_dly0 = '1'
    -----------------------------------------------------------------------------
    TXD_RDY_INDICATOR : process (AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rdy <= '0';
        else
          if clr_txd_rdy = '1' then
            txd_rdy <= '0';
          elsif set_txd_rdy = '1' then
            txd_rdy <= '1';
          else
            txd_rdy <= txd_rdy;
          end if;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Filter to indicate first packet was written
    --    Needed for full flag
    -----------------------------------------------------------------------------
    FIRST_PACKET_WROTE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          wrote_first_packet <= '0';
        elsif set_first_packet = '1' then
          wrote_first_packet <= '1';
        else
          wrote_first_packet <= wrote_first_packet;
        end if;
      end if;
    end process;


    axi_str_txd_2_mem_addr_int_plus1 <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 1);
    axi_str_txd_2_mem_addr_int_plus2 <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 2);
    axi_str_txd_2_mem_addr_int_plus3 <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 3);
    axi_str_txd_2_mem_addr_int_plus4 <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 4);


    ---------------------------------------------------------------------------
    --  Register to help fmax
    --  With ASYNC BRAM clock cannot read/write same address in memory at same
    --  time unless timing is met, so read until data matches
    ---------------------------------------------------------------------------
    RD_PNTR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rd_pntr_1 <= (others => '0');
          txd_rd_pntr   <= (others => '0');
          compare_addr0_cmplt <= '0';
        else
          if set_txc_addr_0 = '1' and txc_addr_0_dly2 = '1' and
             txc_we_dly2 = '0'  then
          --  txc_addr_0_dly2 is when data is first avaliable from memory

          --  use set_txc_addr_0 to disable compare_addr0_cmplt once pointers update
          --  once state machine advances, set_txc_addr_0 will go low so use it to disable any more
          --  any more data from memory
            txd_rd_pntr_1      <= Axi_Str_TxC_2_Mem_Dout(c_TxD_addrb_width -1 downto 0);

            if Axi_Str_TxC_2_Mem_Dout(c_TxD_addrb_width -1 downto 0) = txd_rd_pntr_1 and
              compare_addr0_cmplt = '0' then
              txd_rd_pntr         <= txd_rd_pntr_1;
              if enable_compare_addr0_cmplt = '1' then
                compare_addr0_cmplt <= '1';
              else
                compare_addr0_cmplt <= '0';
              end if;
            else
              txd_rd_pntr         <= txd_rd_pntr;
              compare_addr0_cmplt <= '0';
            end if;
          else
            txd_rd_pntr_1      <= txd_rd_pntr_1;
            txd_rd_pntr        <= txd_rd_pntr;
            compare_addr0_cmplt<= '0';
          end if;
        end if;
      end if;
    end process;


    ---------------------------------------------------------------------------
    --  Update the read pointer locations until the memory goes FULL
    --    Then use the stored values to compare against real time read pointer
    --    and throttle appropriately
    ---------------------------------------------------------------------------
    RD_PNTRS : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rd_pntr_hold_plus3 <= txc_rd_addr3;
          txd_rd_pntr_hold       <= txc_rd_addr0;
        else
          if (txd_mem_full = '0' and txc_addr_0_dly2 = '1' and halt_pntr_update = '0') or update_rd_pntrs = '1'then -- wait on this as it might not be needed  or update_hold_pntrs = '1' then --and
          --  halt_pntr_update is for the special case when memory is almost full/full and
          --  the Txd FSM needs to wait for a few reads before the next packet starts
          --  The TxD FSM will assert it HIGH to prevent the poiners from being updated
            txd_rd_pntr_hold_plus3 <= std_logic_vector(unsigned(txd_rd_pntr) +3);
            txd_rd_pntr_hold       <= txd_rd_pntr;
          else
            txd_rd_pntr_hold_plus3 <= txd_rd_pntr_hold_plus3;
            txd_rd_pntr_hold       <= txd_rd_pntr_hold;
          end if;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Full flag indicator
    --    Does not begin comparison until 1st packet is written to memory
    -----------------------------------------------------------------------------
    TXD_FULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
            txd_mem_full     <= '0';
            txd_mem_not_full <= '1';
        else
            if (axi_str_txd_2_mem_addr_int_plus3 = txd_rd_pntr and
                (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) or
               set_txd_mem_full = '1' then
              txd_mem_full     <= '1';
              txd_mem_not_full <= '0';
            else
              txd_mem_full     <= txd_mem_full;
              txd_mem_not_full <= txd_mem_not_full;
            end if;
        end if;
      end if;
    end process;

    TXD_AFULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
            txd_mem_afull     <= '0';
        else

          if (axi_str_txd_2_mem_addr_int_plus4 = txd_rd_pntr and
              (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) or
             set_txd_mem_afull = '1' then
            txd_mem_afull     <= '1';
          else
            txd_mem_afull     <= txd_mem_afull;
          end if;
        end if;
      end if;
    end process;

    DELAY_TXD_TREADY_DISABLE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        disable_txd_trdy_dly <= disable_txd_trdy;
      end if;
    end process;

    DELAY_TREADY_DISABLE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        disable_txc_trdy_dly <= disable_txc_trdy;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  TxD Ready
    --    Only assert when FIFO is not full and TxC is not in process
    -----------------------------------------------------------------------------
    TXD_READY : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_tready_int_dly <= axi_str_txd_tready_int;
        if (AXI_STR_TXD_TLAST = '1' and AXI_STR_TXD_TVALID = '1' and axi_str_txd_tready_int = '1') or
           (clr_txd_trdy = '1' and disable_txd_trdy_dly = '0') or
           disable_txd_trdy = '1' then
          axi_str_txd_tready_int <= '0';
        elsif set_txd_rdy = '1' or (txd_rdy = '1' and clr_txd_rdy = '0') then
            if (axi_str_txd_2_mem_addr_int_plus3 = txd_rd_pntr and
               inc_txd_wr_addr = '1') or
               (clr_full_pntr = '0' and txd_mem_full = '1') then
            --  txd_rd_pntr is where the the current read is occuring, so
            --    to account for register pipelines, this needs to stop at
            --    3 counts before the current write address
              axi_str_txd_tready_int <= '0';
            else
              axi_str_txd_tready_int <= '1';
            end if;
        else
          axi_str_txd_tready_int <= '0';
        end if;
      end if;
    end process;

    AXI_STR_TXD_TREADY     <= axi_str_txd_tready_int;


    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_WR_ADDR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_2_mem_addr_int       <= (others => '0');
          axi_str_txd_2_mem_addr_int_mins1 <= (others => '0');
        elsif (inc_txd_wr_addr = '1' or inc_txd_addr_one = '1') then
        --  the address ready for the next transaction
          axi_str_txd_2_mem_addr_int       <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 1);
          axi_str_txd_2_mem_addr_int_mins1 <= axi_str_txd_2_mem_addr_int;
        elsif wr_hdr_csum = '1' then
          axi_str_txd_2_mem_addr_int       <= csum_ipv4_hdr_addr;
          axi_str_txd_2_mem_addr_int_mins1 <= axi_str_txd_2_mem_addr_int_mins1;
        elsif ptcl_csum_cmplt = '1' and do_full_csum = '1' then
        -- Set the address for the TCP/UDP csum
          axi_str_txd_2_mem_addr_int       <= csum_ptcl_addr;
          axi_str_txd_2_mem_addr_int_mins1 <= axi_str_txd_2_mem_addr_int_mins1;
        elsif csum_en_dly = '1' then
          axi_str_txd_2_mem_addr_int       <= axi_str_txd_2_mem_addr_int_last;
          axi_str_txd_2_mem_addr_int_mins1 <= axi_str_txd_2_mem_addr_int_mins1;
        else
          axi_str_txd_2_mem_addr_int       <= axi_str_txd_2_mem_addr_int;
          axi_str_txd_2_mem_addr_int_mins1 <= axi_str_txd_2_mem_addr_int_mins1;
        end if;
      end if;
    end process;


    ---------------------------------------------------------------------------
    --  Force and update the BRAM with the axi_str_txd_2_mem_addr_int
    --  every ~128 writes (~512 bytes)
    ---------------------------------------------------------------------------
    BRAM_UPDATE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_txd_rdy = '1' then
          update_bram_cnt     <= (others => '0');
        else
          if update_bram_cnt(7) = '1' and inc_txd_wr_addr = '1' then
            update_bram_cnt <= ('0' & update_bram_cnt(6 downto 0)) + 1;
          elsif inc_txd_wr_addr = '1' then
            update_bram_cnt <= update_bram_cnt + 1;
          else
            update_bram_cnt <= update_bram_cnt;
          end if;
        end if;
      end if;
    end process;



    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_WR_ADDR_LAST : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_2_mem_addr_int_last <= (others => '0');
        elsif wr_hdr_csum = '1' then
        --  hold TxD address to restore after CSUM is written
          axi_str_txd_2_mem_addr_int_last <= axi_str_txd_2_mem_addr_int;
        else
          axi_str_txd_2_mem_addr_int_last <= axi_str_txd_2_mem_addr_int_last;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay the CSUM enable to resore the memory address after the CSUM value
    --  is written
    -----------------------------------------------------------------------------
    CSUM_ENABLE_DELAY : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        -- Used to restore the BRAM Address after writing the Header CSUM and TCP/UDP CSUM
        csum_en_dly <= wr_hdr_csum or (ptcl_csum_cmplt and do_full_csum);    --279 byte sim issue changed do_csum to do_full_csum
      end if;                                                                -- set address back to zero after first packet
    end process;


    axi_str_txd_2_mem_addr               <= axi_str_txd_2_mem_addr_int;


    Axi_Str_TxD_2_Mem_Din(35)           <= axi_str_txd_2_mem_we_int(3);
    Axi_Str_TxD_2_Mem_Din(26)           <= axi_str_txd_2_mem_we_int(2);
    Axi_Str_TxD_2_Mem_Din(17)           <= axi_str_txd_2_mem_we_int(1);
    Axi_Str_TxD_2_Mem_Din(8)            <= axi_str_txd_2_mem_we_int(0);

    Axi_Str_TxD_2_Mem_Din(34 downto 27) <= axi_str_txd_tdata_dly1(31 downto 24);
    Axi_Str_TxD_2_Mem_Din(25 downto 18) <= axi_str_txd_tdata_dly1(23 downto 16);
    Axi_Str_TxD_2_Mem_Din(16 downto  9) <= axi_str_txd_tdata_dly1(15 downto  8);
    Axi_Str_TxD_2_Mem_Din(7  downto  0) <= axi_str_txd_tdata_dly1( 7 downto  0);

    -----------------------------------------------------------------------------
    --  Write Parity bits to the AXI Stream Data Memory
    --    The parity bit always should be the AXI_STR_TXD_TSTRB bits delayed
    --    except when writing the CSUM value.  If writing CSUM, these bits need
    --    set HIGH for the Half word being written; otherwise, the transmission
    --    will end prematurely.
    -----------------------------------------------------------------------------
    MEM_TXD_PARITY : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if wr_hdr_csum = '1' then
          axi_str_txd_2_mem_we_int <= csum_ipv4_hdr_we;
        elsif ptcl_csum_cmplt = '1' and do_full_csum = '1' then
          -- Write the memory with the csum enable bits
          axi_str_txd_2_mem_we_int <= csum_ptcl_we;
        else
          axi_str_txd_2_mem_we_int <= set_txd_we;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Write Enable bits to the AXI Stream Data Memory
    --    All of the write enables bits should be forced HIGH any time a write to
    --    memory is being performed (except csum).  This will allow the parity
    --    bits to be cleared which in turn prevents too much data being read on
    --    the Txd client interface.
    --  When CSUM is being performed, only set the WEs for the half word being
    --  accessed.
    -----------------------------------------------------------------------------
    MEM_TXD_WR_EN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if wr_hdr_csum = '1' then
          Axi_Str_TxD_2_Mem_We <= csum_ipv4_hdr_we;
        elsif ptcl_csum_cmplt = '1' and do_full_csum = '1' then
          -- Set the memory enable bits to allow the CSUM ddata to be written
          Axi_Str_TxD_2_Mem_We <= csum_ptcl_we;
        else
          case set_txd_we is
            when "0000" => Axi_Str_TxD_2_Mem_We <= "0000";
            when others => Axi_Str_TxD_2_Mem_We <= "1111";
          end case;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Enable bit to the AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_EN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if set_txd_en = '1' or wr_hdr_csum = '1' or (ptcl_csum_cmplt = '1' and do_full_csum = '1') then
          -- Enable the memory to be written with the CSUM calculations
          axi_str_txd_2_mem_en_int <= '1';
        else
          axi_str_txd_2_mem_en_int <= '0';
        end if;
      end if;
    end process;

    Axi_Str_TxD_2_Mem_En <= axi_str_txd_2_mem_en_int;

-------------------------------------------------------------------------------
--  End Full CSUM
-------------------------------------------------------------------------------

end rtl;


------------------------------------------------------------------------------
-- tx_vlan_if.vhd
------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- tx_vlan_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_vlan_if.vhd
-- Version:         v1.00a
-- Description:     top level of embedded ip Ethernet MAC interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--                    tx_axistream_if.vhd
--                      tx_basic_if.vhd
--                      tx_csum_if.vhd
--                        tx_csum_partial_if.vhd
--                          tx_csum_partial_calc_if.vhd
--                        tx_full_csum_if.vhd
--          ->          tx_vlan_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tx_if_pack.all;




------------------------------------------------------------------------------
-- Port Declaration
------------------------------------------------------------------------------

entity tx_vlan_if is
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_TYPE                 : integer range 0 to 2         := 0;
    C_PHY_TYPE             : integer range 0 to 7         := 1;
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data

    --Transmit EMAC Interface

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0);  --  Tx AXI-Stream Control to Memory Full Flag

    tx_vlan_bram_addr      : out std_logic_vector(11 downto 0);                     --  Transmit VLAN BRAM Addr
    tx_vlan_bram_din       : in  std_logic_vector(13 downto 0);                     --  Transmit VLAN BRAM Rd Data
    tx_vlan_bram_en        : out std_logic;                                         --  Transmit VLAN BRAM Enable

    enable_newFncEn        : out std_logic; --Only perform VLAN when the FLAG = 0xA --  Enable Extended VLAN Functions
    transMode_cross        : in  std_logic;                                         --  VLAN Translation Mode Control Bit
    tagMode_cross          : in  std_logic_vector( 1 downto 0);                     --  VLAN TAG Mode Control Bits
    strpMode_cross         : in  std_logic_vector( 1 downto 0);                     --  VLAN Strip Mode Control Bits

    tpid0_cross            : in  std_logic_vector(15 downto 0);                     --  VLAN TPID
    tpid1_cross            : in  std_logic_vector(15 downto 0);                     --  VLAN TPID
    tpid2_cross            : in  std_logic_vector(15 downto 0);                     --  VLAN TPID
    tpid3_cross            : in  std_logic_vector(15 downto 0);                     --  VLAN TPID

    newTagData_cross       : in  std_logic_vector(31 downto 0)                      --  VLAN Tag Data

  );
end tx_vlan_if;

architecture rtl of tx_vlan_if is


   --------------------------------------------------------------------------
   -- Signal Declarations
   --------------------------------------------------------------------------
   --Signals for State Machine
   signal set_vlan_bram_en       : std_logic;
   signal clr_vlan_bram_en       : std_logic;
   signal tx_vlan_bram_en_int    : std_logic;
   signal tx_vlan_bram_en_dly1   : std_logic;
   signal tx_vlan_bram_en_dly2   : std_logic;
   
   signal set_decode_dly         : std_logic;
   signal decode_dly1            : std_logic;   
   signal decode_dly2            : std_logic;   
   signal decode_dly3            : std_logic;
   signal decode_dly4            : std_logic;  
   signal inhibit_checktag0tpid  : std_logic;    
   signal tx_vlan_bram_din_dly   : std_logic_vector(13 downto 0);
   signal tx_vlan_bram_addr_int  : std_logic_vector(11 downto 0);



   signal setCheckTag0Tpid       : std_logic;
   signal checkTag0Tpid          : std_logic;
   signal checkTag0Tpid_dly1     : std_logic;
   signal checkTag0Tpid_dly      : std_logic;

   signal setCheckTag1Tpid       : std_logic;
   signal checkTag1Tpid          : std_logic;
   signal checkTag1Tpid_dly1     : std_logic;
   signal checkTag1Tpid_dly      : std_logic;

   signal clr_all_hits             : std_logic;

   --  VLAN Control Signals
   signal tag0TpidHit            : std_logic;
   signal tag0TpidHit_int        : std_logic;
   signal tag1TpidHit            : std_logic;
   signal tag1TpidHit_int        : std_logic;
   signal bramDinTag0Reg         : std_logic;
   signal tag0TpidHitReg         : std_logic;
   signal tag0TotalHit           : std_logic;
   signal newTagTotalHit         : std_logic;
   signal transTotalHit          : std_logic;
   signal transReg               : std_logic_vector(11 downto 0);

  constant zeroes_txc            : std_logic_vector(c_TxC_write_width_b -1 downto c_TxC_addrb_width) := (others => '0');
  constant zeroes_txd            : std_logic_vector(c_TxC_write_width_b -1 downto c_TxD_addrb_width) := (others => '0');
  constant zeroes_txd_2          : std_logic_vector(c_TxC_write_width_b -1 downto c_TxD_addrb_width + 2 ) := (others => '0');

  type TXC_WR_FSM_TYPE is (
                       TXC_ADDR2_WR,
                       TXC_ADDR0_WR,
                       WAIT_WR_CMPLT,
                       TXC_WD0,
--                       WAIT_TXD_FULL,
                       TXC_WD1,
                       WAIT_ADDR2_COMPARE_CMPLT,--added for BRAM async clocks
                       TXC_WD2,
                       TXC_WD3,
                       TXC_WD4,
                       WAIT_ADDR0_COMPARE_CMPLT,--added for BRAM async clocks
                       TXC_WD5,
                       WAIT_TXD_CMPLT,
                       WAIT_TXD_MEM,
                       WR_TXC_PNTR,
                       WR_TXD_END_PNTR
                      );
  signal txc_wr_cs, txc_wr_ns             : TXC_WR_FSM_TYPE;

  type TXD_WR_FSM_TYPE is (
                       IDLE,
                       DST_SRC,
                       SRC,
                       VLAN1,
                       WAIT_TVALID,
                       VLAN2,
                       DECODE,
                       STTr,
                       STRIP,
                       TAG,
                       TRANSLATE,
                       WAIT_STATE,
                       TXD_PRM,
                       TXD_WRT,
                       MEM_FULL,
                       CLR_WORDS,
                       WAIT_WR1,
                       WAIT_WR2,
                       WAIT_COMPARE_CMPLT
                      );
  signal txd_wr_cs, txd_wr_ns             : TXD_WR_FSM_TYPE;

  signal txc_min_wr_addr                  : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_rsvd_wr_addr                 : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_max_wr_addr                  : std_logic_vector(c_TxC_addrb_width -1 downto 0);

  signal txc_wr_addr0                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr1                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr2                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr3                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr5                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr6                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);

  signal axi_str_txc_tready_int           : std_logic;
  signal axi_str_txc_tready_int_dly       : std_logic;
  signal axi_str_txc_tvalid_dly0          : std_logic;
  signal axi_str_txc_tlast_dly0           : std_logic;
--  signal axi_str_txc_tstrb_dly0           : std_logic_vector(3 downto 0);
  signal axi_str_txc_tdata_dly0           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal clr_txc_trdy                     : std_logic;

  signal axi_str_txd_tready_int           : std_logic;
  signal axi_str_txd_tready_int_dly       : std_logic;
  signal axi_str_txd_tvalid_dly0          : std_logic;
  signal axi_str_txd_tlast_dly0           : std_logic;
  signal axi_str_txd_tstrb_dly0           : std_logic_vector(3 downto 0);
  signal axi_str_txd_tdata_dly0           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal axi_str_txd_tdata_dly1           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal clr_txd_trdy                     : std_logic;

  signal set_txc_addr_0                   : std_logic;
  signal txc_addr_0_dly1                  : std_logic;
  signal txc_addr_0_dly2                  : std_logic;
  signal set_txc_addr_1                   : std_logic;
  signal txc_addr_1                       : std_logic;
  signal set_txc_addr_2                   : std_logic;
  signal txc_addr_2                       : std_logic;
  signal set_txc_addr_4_n                 : std_logic;
  signal set_txc_addr_3                   : std_logic;
  signal clr_txc_addr_3                   : std_logic;
  signal txc_addr_3_dly                   : std_logic;
  signal txc_addr_3_dly2                  : std_logic;
  signal txc_addr_3_dly3                  : std_logic;
  signal inc_txd_addr_one                 : std_logic;
  signal set_txc_trdy                     : std_logic;
  signal set_txc_trdy2                    : std_logic;
  signal clr_txc_trdy2                    : std_logic;
  signal set_txcwr_rd_addr                : std_logic;
  signal set_txcwr_wr_end                 : std_logic;
  signal set_txc_en                       : std_logic;
  signal set_txc_we                       : std_logic;
  signal txc_we                           : std_logic;
  signal txc_we_dly1                      : std_logic;
  signal txc_we_dly2                      : std_logic;
  signal addr_2_en                        : std_logic;
  signal addr_2_en_dly1                   : std_logic;
  signal addr_2_en_dly2                   : std_logic;

  signal txc_mem_full                     : std_logic;
  signal txc_mem_not_full                 : std_logic;
  signal txc_mem_afull                    : std_logic;
  signal txc_mem_wr_addr                  : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_0                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_1                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_last             : std_logic_vector(c_TxC_addrb_width   -1 downto 0);

  signal Axi_Str_TxC_2_Mem_Addr_int       : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal Axi_Str_TxC_2_Mem_We_int         : std_logic_vector(0 downto 0);
  signal txc_mem_wr_addr_plus1            : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_plus2            : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_rd_addr2_pntr                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_rd_addr2_pntr_1              : std_logic_vector(c_TxC_addrb_width   -1 downto 0);


  -- Set to the full width of the write data bus
  signal Axi_Str_TxC_2_Mem_Din_int        : std_logic_vector(c_TxC_write_width_b -1 downto 0);

  signal set_axi_flag                     : std_logic;
  signal set_csum_cntrl                   : std_logic;
  signal set_csum_begin_insert            : std_logic;
  signal set_csum_rsvd_init               : std_logic;
  signal axi_flag                         : std_logic_vector( 3 downto 0);
  signal csum_cntrl                       : std_logic_vector( 1 downto 0);

  signal set_first_packet                 : std_logic;
  signal wrote_first_packet               : std_logic;
  signal inc_txd_wr_addr                  : std_logic;
  signal set_txd_we                       : std_logic_vector( 3 downto 0);
  signal set_txd_en                       : std_logic;
  signal set_txd_rdy                      : std_logic;
  signal clr_txd_rdy                      : std_logic;
  signal clr_full_pntr                    : std_logic;
  signal halt_pntr_update                 : std_logic;
  signal disable_txd_trdy                 : std_logic;
  signal disable_txd_trdy_dly             : std_logic;
  signal disable_txc_trdy                 : std_logic;
  signal disable_txc_trdy_dly             : std_logic;

  signal txd_rdy                          : std_logic;
  signal axi_str_txd_2_mem_addr_int       : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus1 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus3 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus4 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus10: std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txd_mem_clr_words                : std_logic;
  signal txd_mem_full                     : std_logic;
  signal txd_mem_not_full                 : std_logic;
  signal txd_mem_afull                    : std_logic;
  signal axi_str_txd_2_mem_we_int         : std_logic_vector( 3 downto 0);
  signal axi_str_txd_2_mem_en_int         : std_logic;

  signal txd_rd_pntr                      : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_1                    : std_logic_vector(c_TxD_addrb_width -1 downto 0);

  signal nine                             : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal update_cnt                       : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_max_wr_addr                  : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_max_wr_addr_minus4           : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_max_wr_addr_minus10          : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_hold_plus3           : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_hold_plus9           : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_hold                 : std_logic_vector(c_TxD_addrb_width -1 downto 0);

  signal vlan_sel                         : std_logic_vector(2 downto 0);
  signal set_mux_dly                      : std_logic;
  signal clr_mux_dly                      : std_logic;
  signal txd_throttle                     : std_logic;
  signal txd_throttle_dly                 : std_logic;
  signal ignore_tvalid                    : std_logic;
  signal ignore_tvalid_dly                : std_logic;
  signal set_txd_tlast_rcvd               : std_logic;
  signal free_up_memory                   : std_logic;
  signal set_mux_tag                      : std_logic;
  signal set_mux_trans                    : std_logic;

  --implement logic below

  signal load_data_1                      : std_logic;
  signal load_data_1_dly                  : std_logic;
  signal set_mux_data_1_reg               : std_logic;
  signal set_mux_tlast_1_reg              : std_logic;

  signal load_data_2                      : std_logic;
  signal set_mux_data_2_reg               : std_logic;
  signal set_mux_tlast_2_reg              : std_logic;

  signal axi_str_txd_tstrb_1              : std_logic_vector(3 downto 0);
  signal axi_str_txd_tstrb_2              : std_logic_vector(3 downto 0);
  signal axi_str_txd_tlast_1              : std_logic;
  signal axi_str_txd_tlast_2              : std_logic;
  signal axi_str_txd_data_1               : std_logic_vector(31 downto 0);
  signal axi_str_txd_data_2               : std_logic_vector(31 downto 0);

  signal ignore_txd_trdy                  : std_logic;
  signal tx_init_in_prog_int              : std_logic;
  signal init_bram                        : std_logic;

  signal txc_rd_addr0                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txc_rd_addr2                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txc_rd_addr3                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txc_rd_addr9                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);

  signal compare_addr0                    : std_logic;
  signal compare_addr0_cmplt              : std_logic;

  signal compare_addr2                    : std_logic;
  signal compare_addr2_cmplt              : std_logic;
  signal compare_addr2_cmplt_dly          : std_logic;

  signal update_bram_cnt                  : std_logic_vector(7 downto 0);

  signal enable_compare_addr0_cmplt       : std_logic;
  signal set_ignore_txd_tvalid            : std_logic;
  signal ignore_txd_tvalid                : std_logic;

  signal end_addr_byte_offset             : std_logic_vector(1 downto 0);
  signal check_full                       : std_logic;
  signal update_rd_pntrs                  : std_logic;
  signal update_rd_pntrs_reg              : std_logic;
  signal first_packet                     : std_logic;
  
  signal set_tag_en_go                    : std_logic; 
  signal tag_en_go                        : std_logic;
  
  
  begin





   --************************************************************************--
   ----------------------------------------------------------------------------
   -- START
   -- -  Strip, Tag, and Translation Hit Logic based upon parameter settings
   --    and register settings
   --
   ----------------------------------------------------------------------------
   ----------------------------------------------------------------------------
   -- Set strip TPID hit if stripping is enabled
   ----------------------------------------------------------------------------
   GEN_TAG0_HIT : if C_TXVLAN_STRP = 1 generate
   begin

      -------------------------------------------------------------------------
      -- Stage 1
      -- Compare delayed TPID value from LLink against the 4 TPID values
      -- stored in SW accessable registers -
      -------------------------------------------------------------------------

      CHECK_TAG0_TPID_HIT : process(AXI_STR_TXD_ACLK)
      begin

        if rising_edge(AXI_STR_TXD_ACLK) then
          if checkTag0Tpid = '1' and inhibit_checktag0tpid = '0' then
            if axi_str_txd_tdata_dly0(15 downto 0) = tpid0_cross(7 downto 0) & tpid0_cross(15 downto 8) or
               axi_str_txd_tdata_dly0(15 downto 0) = tpid1_cross(7 downto 0) & tpid1_cross(15 downto 8) or
               axi_str_txd_tdata_dly0(15 downto 0) = tpid2_cross(7 downto 0) & tpid2_cross(15 downto 8) or
               axi_str_txd_tdata_dly0(15 downto 0) = tpid3_cross(7 downto 0) & tpid3_cross(15 downto 8) then
               tag0TpidHit_int <= '1';
            else
               tag0TpidHit_int <= '0';
            end if;
          else
            tag0TpidHit_int <= '0';
          end if;

          tag0TpidHit <= tag0TpidHit_int;

        end if;
      end process;


      ----------------------------------------------------------------------------
      -- This process is needed to hold the BRAM Data and tag0 hit data until a
      -- decision can be made on which data to translate
      -- - data from this read or data from the next read
      --  - the last clock cycle tx_vlan_bram_en_dly1 is HIGH will capture the
      --    BRAM TAG bit from the first VLAN TAG
      ----------------------------------------------------------------------------
      REG_BRAM_DOUT_A_TAG_0 : process(AXI_STR_TXD_ACLK)
      begin

         if rising_edge(AXI_STR_TXD_ACLK) then
            if reset2axi_str_txd = '1' or clr_all_hits = '1' then
               bramDinTag0Reg <= '0';
--            elsif checkTag0Tpid_dly = '1' then
            elsif checkTag0Tpid_dly = '1' then
               bramDinTag0Reg <= tx_vlan_bram_din_dly(0);
            else
               bramDinTag0Reg <= bramDinTag0Reg;
            end if;
         end if;
      end process;


      ----------------------------------------------------------------------------
      -- If the TPID from tag0 is a hit then save this data in case a
      -- strip does not occure.  Then if a tag occurs, the data will be available
      ----------------------------------------------------------------------------
      REG_TAG0_TPID_HIT : process(AXI_STR_TXD_ACLK)
      begin

         if rising_edge(AXI_STR_TXD_ACLK) then
            if reset2axi_str_txd = '1' or clr_all_hits = '1' then
               tag0TpidHitReg   <= '0';
            elsif tag0TpidHit = '1' then
               tag0TpidHitReg   <= '1';
            elsif axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
               tag0TpidHitReg   <= '0';
            else
               tag0TpidHitReg <= tag0TpidHitReg;
            end if;
         end if;
      end process;


      ----------------------------------------------------------------------------
      -- Stage 2
      -- If tag0TotalHit is set, then check the strip mode bits to determine
      -- how/if a total hit occurs.
      --    If strpMode_cross = 00 then no stripping occures
      --    If strpMode_cross = 01 then only strip if it is a VLAN tag
      --       ie if tag0TotalHit=1
      --    If strpMode_cross = 10 then do not strip anything
      --       this mode is reserved and has no function
      --    If strpMode_cross = 11 then strip select VLAN frames based upon:
      --       1. Must be a VLAN Hit (tag0TotalHit must be set) and
      --       2. tx_vlan_bram_din_dly Strip Enable bit must be set
      ----------------------------------------------------------------------------
      SET_TAG0_HIT : process(AXI_STR_TXD_ACLK)
      begin

         if rising_edge(AXI_STR_TXD_ACLK) then
            if reset2axi_str_txd = '1' or clr_all_hits = '1' then
               tag0TotalHit <= '0';
            else
               case strpMode_cross is
                  when "11"   =>
                  -- Strip one tag from select VLAN tagged frames
                     if tag0TpidHit = '1' then
                        tag0TotalHit <= tx_vlan_bram_din_dly(1);
                     else
                        tag0TotalHit <= tag0TotalHit;
                     end if;
                  when "01"   =>
                  -- Strip one tagg from all VLAN tagged frames
                     if tag0TpidHit = '1' then
                        tag0TotalHit <= '1';
                     else
                        tag0TotalHit <= tag0TotalHit;
                     end if;
                  when others =>
                  -- do not strip any tags
                     tag0TotalHit <= '0';
               end case;
            end if;
         end if;
      end process;

   end generate;


   ----------------------------------------------------------------------------
   -- Stage 1 and Stage 2
   -- Force strip hit low when stripping is not enabled
   ----------------------------------------------------------------------------
   GEN_NO_TAG0_HIT : if C_TXVLAN_STRP = 0 generate
   begin

      tag0TotalHit   <= '0';
      tag0TpidHit    <= '0';
      tag0TpidHit_int<= '0';
      tag0TpidHitReg <= '0';
      bramDinTag0Reg <= '0';
   end generate;



   ----------------------------------------------------------------------------
   -- Stage 1
   -- Compare delayed TPID value from LLink against the 4 TPID values stored in
   -- SW accessable registers -
   -- -  Without stripping enabled checkTag0Tpid occurs on the 4th 32-bit LL
   --    Data word (the first word after the SRC Address)
   ----------------------------------------------------------------------------
   GEN_TRANS_TAG_HIT_NO_STRIP : if ((C_TXVLAN_TRAN = 1 or C_TXVLAN_TAG = 1) and
                                     C_TXVLAN_STRP = 0) generate
   begin


      CHECK_TRANS_TAG_TPID_HIT : process(AXI_STR_TXD_ACLK)
      begin

        if rising_edge(AXI_STR_TXD_ACLK) then
          if checkTag0Tpid = '1' and inhibit_checktag0tpid = '0' then
            if axi_str_txd_tdata_dly0(15 downto 0) = tpid0_cross(7 downto 0) & tpid0_cross(15 downto 8) or
               axi_str_txd_tdata_dly0(15 downto 0) = tpid1_cross(7 downto 0) & tpid1_cross(15 downto 8) or
               axi_str_txd_tdata_dly0(15 downto 0) = tpid2_cross(7 downto 0) & tpid2_cross(15 downto 8) or
               axi_str_txd_tdata_dly0(15 downto 0) = tpid3_cross(7 downto 0) & tpid3_cross(15 downto 8) then
               tag1TpidHit_int <= '1';
            else
               tag1TpidHit_int <= '0';
            end if;
          else
            tag1TpidHit_int <= '0';
          end if;

          tag1TpidHit <= tag1TpidHit_int;

        end if;
      end process;
   end generate;


   ----------------------------------------------------------------------------
   -- Stage 1
   -- Compare delayed TPID value from LLink against the 4 TPID values stored in
   -- SW accessable registers -
   -- -  With stripping enabled checkTag1Tpid occurs on the 5th 32-bit LL Data
   --    word (the second word after the SRC Address)
   ----------------------------------------------------------------------------
   GEN_TRANS_TAG_HIT_WITH_STRIP : if ((C_TXVLAN_TRAN = 1 or C_TXVLAN_TAG = 1) and
                                       C_TXVLAN_STRP = 1) generate
   begin



      CHECK_TRANS_TAG_TPID_HIT : process(AXI_STR_TXD_ACLK)
      begin

        if rising_edge(AXI_STR_TXD_ACLK) then
          if checkTag1Tpid = '1' and axi_str_txd_tvalid_dly0 = '1' then
          --  axi_str_txd_tdata can change while tvalid is low, so do not allow compare until
          --  axi_str_txd_tvalid_dly0 is HIGH
            if axi_str_txd_tdata_dly0(15 downto 0) = tpid0_cross(7 downto 0) & tpid0_cross(15 downto 8) or
               axi_str_txd_tdata_dly0(15 downto 0) = tpid1_cross(7 downto 0) & tpid1_cross(15 downto 8) or
               axi_str_txd_tdata_dly0(15 downto 0) = tpid2_cross(7 downto 0) & tpid2_cross(15 downto 8) or
               axi_str_txd_tdata_dly0(15 downto 0) = tpid3_cross(7 downto 0) & tpid3_cross(15 downto 8) then
               tag1TpidHit_int <= '1';
            else
               tag1TpidHit_int <= '0';
            end if;
          else
            tag1TpidHit_int <= '0';
          end if;

          tag1TpidHit <= tag1TpidHit_int;

        end if;
      end process;
   end generate;


   ----------------------------------------------------------------------------
   -- Stage 1
   -- Compare delayed TPID value from LLink against the 4 TPID values stored in
   -- SW accessable registers -
   ----------------------------------------------------------------------------
   GEN_NO_TRANS_TAG_HIT : if (C_TXVLAN_TRAN = 0 and C_TXVLAN_TAG = 0) generate
   begin

      tag1TpidHit <= '0';
   end generate;


   ----------------------------------------------------------------------------
   -- Stage 2
   -- Set tag total hit only if tagging is enabled and the mode allows it
   --    If  tagMode_cross = "00" then do NOT tag any frames
   --    If  tagMode_cross = "01" then tag all frames even if it was not a
   --       VLAN HIT (tag1TpidHit = '0')
   --    If  tagMode_cross = "10" then add one tag to all VLAN Frames
   --       (tag1TpidHit = '1')
   --    If  tagMode_cross = "11" then add one tag to select VLAN frames
   --       based upon the tx_vlan_bram_din_dly tag bit being set
   --
   --       HOWEVER, since stripping is enabled, must decide which TAG to
   --       evaluate for  setting newTagTotalHit
   --          If a strip is occuring, then use the inner TAG
   --          If a strip is not going to occur, use the outer TAG
   ----------------------------------------------------------------------------
   GEN_TAG_HIT_WITH_STRIP : if C_TXVLAN_TAG = 1 and C_TXVLAN_STRP = 1 generate
   begin

      SET_TAG_HIT : process(AXI_STR_TXD_ACLK)
      begin

         if rising_edge(AXI_STR_TXD_ACLK) then
            if reset2axi_str_txd = '1' or clr_all_hits = '1' then
               newTagTotalHit <= '0';
            else
               case tagMode_cross is
                  when "11"   =>
                  --  Only tag select VLAN tagged frames
                     -- Strip is going to occur, so newTagTotalHit is set
                     -- by tpid hit from 2nd tag (tag1TpidHit)
                     if tag0TotalHit = '1' then
                        if tag1TpidHit = '1' then
                           newTagTotalHit <= tx_vlan_bram_din_dly(0);
                        else
                           newTagTotalHit <= newTagTotalHit;
                        end if;
                     else
                     -- Otherwise a strip is not occuring, so newTagTotalHit is
                     -- set by the tpid from the previous tag (tag0TpidHitReg)
                        if tag0TpidHitReg = '1' then
                           newTagTotalHit <= bramDinTag0Reg;
                        else
                           newTagTotalHit <= newTagTotalHit;
                        end if;
                     end if;

                  when "10"   =>
                  --  Only tag VLAN tagged frames
                     -- Strip is going to occur, so newTagTotalHit is set
                     -- by tpid hit from 2nd tag (tag1TpidHit)
                     if tag0TotalHit = '1' then  --strip will occur
                        if tag1TpidHit = '1' then  --2nd Tag hit
                           newTagTotalHit <= '1';
                        else
                           newTagTotalHit <= newTagTotalHit;
                        end if;
                     else
                     -- Otherwise a strip is not occuring, so newTagTotalHit is
                     -- set by the tpid from the previous tag (tag0TpidHitReg)
                        if tag0TpidHitReg = '1' then
                           newTagTotalHit <= '1';
                        else
                           newTagTotalHit <= newTagTotalHit;
                        end if;
                     end if;
                  when "01"   =>
                  --  Tag ALL frames
                     if checkTag1Tpid_dly = '1' then
                        newTagTotalHit <= '1';
                     else
                        newTagTotalHit <= newTagTotalHit;
                     end if;
                  when others =>
                  --  Do not tag any frames
                     newTagTotalHit <= '0';
               end case;
            end if;
         end if;
      end process;

   end generate;


   ----------------------------------------------------------------------------
   -- Stage 2
   -- Set tag total hit only if tagging is enabled and the mode allows it
   --    If  tagMode_cross = "00" then do NOT tag any frames
   --    If  tagMode_cross = "01" then tag all frames even if it was not a
   --       VLAN HIT (tag1TpidHit = '0')
   --    If  tagMode_cross = "10" then add one tag to all VLAN Frames
   --       (tag1TpidHit = '1')
   --    If  tagMode_cross = "11" then add one tag to select VLAN frames
   --       based upon the tx_vlan_bram_din_dly tag bit being set
   --
   --    Always use the outer TAG when stripping is disabled by the parameter
   ----------------------------------------------------------------------------
   GEN_TAG_HIT_NO_STRIP : if C_TXVLAN_TAG = 1 and C_TXVLAN_STRP = 0 generate
   begin

      SET_TAG_HIT : process(AXI_STR_TXD_ACLK)
      begin

         if rising_edge(AXI_STR_TXD_ACLK) then
            if reset2axi_str_txd = '1' or clr_all_hits = '1' then
               newTagTotalHit <= '0';
            else
               case tagMode_cross is
                  when "11"   =>
                  --  Only tag select VLAN tagged frames
                     if tag1TpidHit = '1' then
                        newTagTotalHit <= tx_vlan_bram_din_dly(0);
                     else
                        newTagTotalHit <= newTagTotalHit;
                     end if;
                  when "10"   =>
                  --  Only tag VLAN tagged frames
                     if tag1TpidHit = '1' then
                        newTagTotalHit <= '1';
                     else
                        newTagTotalHit <= newTagTotalHit;
                     end if;
                  when "01"   =>
                  --  Tag ALL frames
                     if checkTag1Tpid_dly = '1' then
                        newTagTotalHit <= '1';
                     else
                        newTagTotalHit <= newTagTotalHit;
                     end if;
                  when others =>
                  --  Do not tag any frames
                     newTagTotalHit <= '0';
               end case;
            end if;
         end if;
      end process;

   end generate;


   ----------------------------------------------------------------------------
   -- Force tag total hit LOW if tagging is NOT enabled
   ----------------------------------------------------------------------------
   GEN_NO_TAG_HIT : if C_TXVLAN_TAG = 0 generate
   begin

      newTagTotalHit <= '0';

   end generate;


   ----------------------------------------------------------------------------
   -- Set translation total hit if translation is enabled
   -- A translation will occure only if transMode_cross is set and a TPID hit occurs
   -- on the first vlan tag when a strip does not occur or the 2nd vlan tag
   -- when a strip does occur.
   ----------------------------------------------------------------------------
   GEN_TRANS_HIT_WITH_STRIP : if C_TXVLAN_TRAN = 1  and C_TXVLAN_STRP = 1 generate
   begin

      SET_TRANS_HIT : process(AXI_STR_TXD_ACLK)
      begin

         if rising_edge(AXI_STR_TXD_ACLK) then
            if reset2axi_str_txd = '1' or clr_all_hits = '1' or transMode_cross = '0' then
               transTotalHit <= '0';
            else
               if tag0TotalHit = '1' then
                  -- Strip is going to occur, so transTotalHit is set
                  -- by tpid hit from 2nd tag (tag1TpidHit)
                  if tag1TpidHit = '1' then
                     transTotalHit <= '1';
                  else
                     transTotalHit <= transTotalHit;
                  end if;
               else
                  -- Otherwise a strip is not occuring, so transTotalHit is
                  -- set by the tpid from the previous tag (tag0TpidHitReg)
                  if tag0TpidHitReg = '1' then
                     transTotalHit <= '1';
                  else
                     transTotalHit <= transTotalHit;
                  end if;
               end if;
            end if;
         end if;
      end process;

   end generate;


   ----------------------------------------------------------------------------
   -- Set translation total hit if translation is enabled
   -- A translation will occure only if transMode_cross is set and a TPID hit occurs
   -- on the first vlan tag since stripping is not enabled.
   ----------------------------------------------------------------------------
   GEN_TRANS_HIT_NO_STRIP : if C_TXVLAN_TRAN = 1  and C_TXVLAN_STRP = 0 generate
   begin

      SET_TRANS_HIT : process(AXI_STR_TXD_ACLK)
      begin

         if rising_edge(AXI_STR_TXD_ACLK) then
            if reset2axi_str_txd = '1' or clr_all_hits = '1' or transMode_cross = '0' then
               transTotalHit <= '0';
            else
               if tag1TpidHit = '1' then
                  transTotalHit <= '1';
               else
                  transTotalHit <= transTotalHit;
               end if;
            end if;
         end if;
      end process;

   end generate;


   ----------------------------------------------------------------------------
   -- Force translate total hit LOW if translation is NOT enabled
   ----------------------------------------------------------------------------
   GEN_NO_TRANS_HIT : if C_TXVLAN_TRAN = 0 generate
   begin

      transTotalHit <= '0';

   end generate;

   ----------------------------------------------------------------------------
   -- Set translation register if translation and stripping parameters are set
   --    It will always load the translation value from the first Bram Read,
   --    then update it with the 2nd Bram read if needed
   --       In either case the loaded data may/may not be used depending upon
   --       if a translation hit occurs
   ----------------------------------------------------------------------------
   GEN_TRANS_REG_WITH_STRIP : if C_TXVLAN_TRAN = 1 and C_TXVLAN_STRP = 1 generate
   begin

      LOAD_TRANS_REG : process(AXI_STR_TXD_ACLK)
      begin

         if rising_edge(AXI_STR_TXD_ACLK) then
            if reset2axi_str_txd = '1' or clr_all_hits = '1' then
               transReg <= (others => '0');
            else
               if checkTag0Tpid_dly = '1' then
               -- Load the first tag into the trans reg
               -- -  This needs to be loaded because the strip may/may not occur at this point
               --    so load it to be safe then check if strip occurs on the next clock
               --    (the condition below)
                  transReg <= tx_vlan_bram_din_dly(13 downto 2);
               elsif tag0TotalHit = '1' and checkTag1Tpid_dly = '1' then
               -- Load the second tag into the trans reg
               -- -  This needs loaded because the first tag is stripped so the
               --    next tag (this one) will be translated
                  transReg <= tx_vlan_bram_din_dly(13 downto 2);
               else
                  transReg <= transReg;
               end if;
            end if;
         end if;
      end process;
   end generate;


   ----------------------------------------------------------------------------
   -- Set translation register if translation aparameter is set
   --    The loaded data may/may not be used depending upon
   --    if a translation hit occurs
   ----------------------------------------------------------------------------
   GEN_TRANS_REG_NO_STRIP : if C_TXVLAN_TRAN = 1 and C_TXVLAN_STRP = 0 generate
   begin

      LOAD_TRANS_REG : process(AXI_STR_TXD_ACLK)
      begin

         if rising_edge(AXI_STR_TXD_ACLK) then
            if reset2axi_str_txd = '1' or clr_all_hits = '1' then
               transReg <= (others => '0');
            else
               if checkTag0Tpid_dly = '1' then
               -- Load the first tag into the trans reg
               -- -  since stripping is not enabled, this is the only tag it can be
                  transReg <= tx_vlan_bram_din_dly(13 downto 2);
               else
                  transReg <= transReg;
               end if;
            end if;
         end if;
      end process;
   end generate;

   ----------------------------------------------------------------------------
   -- Translation is disabled
   ----------------------------------------------------------------------------
   GEN_NO_TRANS_REG : if C_TXVLAN_TRAN = 0 generate
   begin

      transReg <= (others => '0');
   end generate;

   ----------------------------------------------------------------------------
   -- Translation and Tagging are disabled
   ----------------------------------------------------------------------------
   GEN_NO_TT_HIT : if C_TXVLAN_TAG = 0 and C_TXVLAN_TRAN = 0 generate
   begin

      newTagTotalHit   <= '0';
      transTotalHit <= '0';
      transReg     <= (others => '0');
   end generate;

   ----------------------------------------------------------------------------
   -- END
   -- -  Strip, Tag, and Translation Hit Logic based upon parameter settings
   --    and register settings
   ----------------------------------------------------------------------------




   ----------------------------------------------------------------------------
   -- This state machine controls the reading/evaluation of data read from
   -- the BRAM and controls all of the muxing of the pipeline to perform
   -- all of the transmit VLAN functions.
   -- It assumes all three VLAN functions are enabled and
   -- branches accordingly based upon register mode settings for stripping and
   -- tagging.
   -- -  Stripping
   --    -  If strpMode_cross = 00 then no stripping occures
   --    -  If strpMode_cross = 01 then only strip if it is a VLAN tag
   --       ie if tag0TotalHit=1
   --    -  If strpMode_cross = 10 then do not strip anything
   --       this mode is reserved and has no function
   --    -  If strpMode_cross = 11 then strip select VLAN frames based upon:
   --       -  1. Must be a VLAN Hit (tag0TotalHit must be set) and
   --       -  2. tx_vlan_bram_din_dly Strip Enable bit must be set
   --
   -- -  Tagging
   --    -  If  tagMode_cross = "00" then do NOT tag any frames
   --    -  If  tagMode_cross = "01" then tag all frames even if it was not a
   --       VLAN HIT (tag1TpidHit = '0')
   --    -  If  tagMode_cross = "10" then add one tag to all VLAN Frames
   --       (tag1TpidHit = '1')
   --    -  If  tagMode_cross = "11" then add one tag to select VLAN frames
   --       based upon the tx_vlan_bram_din_dly tag bit being set
   --
   -- -  Translation
   --    -  If C_TXVLAN_TRAN is set and the current packet is a VLAN
   --       packet (transTotalHit gets set HIGH), a translation will occur
   --
   -- The state machine transitions from state to state dependant upon
   -- axi_str_txd_tvalid_dly0 and axi_str_txd_tready_int_dly both being LOW, or
   -- if payLoadSizes1_14 is set.  Depending upon the branch taken for VLAN
   -- support, the state machine will stall without this signal for packet
   -- sizes less than 15 (T/L = 0xF).
   ----------------------------------------------------------------------------

    -----------------------------------------------------------------------------
    --  The TxC BRAM is set up to to always store the current TxD Read and Write
    --    pointers in the first two locations (0x0 and 0x1) of the Memory
    --    respectivively.  The current TxC Read and write pointer are always
    --    stored in the the next two locations (0x2 and 0x3) of the Memory
    --    respectively.  The End addresses for each packet are then stored
    --    in the remaing Memory locations starting at address 0x4.  After
    --    the end pointer to the maximum address has been written, if the
    --    memory is not full, the address pointer will loop back to address
    --    0x4 and write the end pointer for the next packet.
    --
    --                                   BRAM
    --                             Write       Read
    --                           _____________________
    --                          |__________|_________| <-- TxD Rd Pointer
    --      TxD Wr Pointer -->  |__________|_________|
    --                          |__________|_________| <-- TxC Rd Pointer
    --      TxC Wr Pointer -->  |__________|_________|
    --      Packet 0 End   -->  |__________|_________|  --> Packet 0 End
    --      Packet 1 End   -->  |__________|_________|  --> Packet 1 End
    --      Packet 2 End   -->  |__________|_________|  --> Packet 2 End
    --         .                |__________|_________|         .
    --         .                |__________|_________|         .
    --         .                |__________|_________|         .
    --      Packet n End   -->  |__________|_________|  --> Packet n End
    --
    -----------------------------------------------------------------------------

    -----------------------------------------------------------------------------
    --  Create the full and empty comparison values for the S6 and V6 since
    --  1 S6 BRAM = 1/2 V6 BRAM
    -----------------------------------------------------------------------------
    GEN_TXC_MIN_MAX_WR_FLAG : for i in (c_TxC_addrb_width-1) downto 0 generate
      txc_min_wr_addr(i)  <= '1' when (i = 2)          else '0'; -- do not loop back to 0x0; loop to 0x4
      txc_max_wr_addr(i)  <= '0' when (i = 0 or i = 1) else '1';
      txc_wr_addr0(i)     <= '0';
      txc_wr_addr1(i)     <= '1' when (i = 0)          else '0';
      txc_wr_addr2(i)     <= '1' when (i = 1)          else '0';
      txc_wr_addr3(i)     <= '1' when (i = 0 or i = 1) else '0';
      txc_wr_addr5(i)     <= '1' when (i = 0 or i = 2) else '0';
      txc_wr_addr6(i)     <= '1' when (i = 1 or i = 2) else '0';
    end generate GEN_TXC_MIN_MAX_WR_FLAG;

    GEN_TXD_MIN_MAX_WR_FLAG : for i in (c_TxD_addrb_width-1) downto 0 generate
      nine(i)                    <= '1' when (i = 0 or i = 3) else '0';
      txd_max_wr_addr_minus4(i)  <= '0' when (i = 2) else '1';
      txd_max_wr_addr_minus10(i) <= '0' when (i = 1 or i = 3) else '1';
      txd_max_wr_addr(i)         <= '1';

    end generate GEN_TXD_MIN_MAX_WR_FLAG;

    GEN_TXC_RD_FLAG : for i in (c_TxD_addrb_width-1) downto 0 generate
      txc_rd_addr0(i)     <= '0';
      txc_rd_addr2(i)     <= '1' when (i = 1)          else '0';
      txc_rd_addr3(i)     <= '1' when (i = 0 or i = 1) else '0';
      txc_rd_addr9(i)     <= '1' when (i = 0 or i = 3) else '0';
    end generate GEN_TXC_RD_FLAG;




    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Control Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXC_CONTROL : process(AXI_STR_TXC_ACLK)
    begin
      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          axi_str_txc_tvalid_dly0 <= '0';
          axi_str_txc_tlast_dly0  <= '0';
          clr_txc_trdy           <= '0';
        else
          axi_str_txc_tvalid_dly0 <= axi_str_txc_tvalid;
          axi_str_txc_tlast_dly0  <= axi_str_txc_tlast;
          if axi_str_txc_tvalid = '1' and axi_str_txc_tlast = '1' and axi_str_txc_tready_int = '1' then
            clr_txc_trdy <= '1';
          else
            clr_txc_trdy <= '0';
          end if;
        end if;
      end if;
    end process;

    -- Register the incoming AXI Stream Control Data Bus
    -----------------------------------------------------------------------------
    REG_TXC_IN : process(AXI_STR_TXC_ACLK)
    begin
      if rising_edge(AXI_STR_TXC_ACLK) then
--          axi_str_txc_tstrb_dly0  <= axi_str_txc_tstrb;
          axi_str_txc_tdata_dly0  <= axi_str_txc_tdata;
      end if;
    end process;    
    
    -----------------------------------------------------------------------------
    --  AXI Stream TX Control State Machine - combinational/combinatorial
    --    Used to register the incoming control and checksum information
    --    This state machine will throttle the Transmit AXI Stream Data state
    --      machine until after the control information has been received.
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXC_CMB : process (txc_wr_cs,axi_str_txc_tvalid_dly0,
      axi_str_txc_tlast_dly0,axi_str_txd_tlast_dly0,
      axi_str_txd_tvalid_dly0,txc_addr_3_dly,
      wrote_first_packet,axi_str_txc_tready_int_dly,axi_str_txd_tready_int_dly,
      disable_txd_trdy_dly,disable_txc_trdy_dly,axi_str_txd_tlast_1,axi_str_txd_tlast_2,
      compare_addr2_cmplt,compare_addr2_cmplt_dly,compare_addr0_cmplt,
      update_bram_cnt,txc_mem_full,load_data_1_dly,tagmode_cross,tag_en_go)
      
    begin


      set_axi_flag               <= '0';
      set_csum_cntrl             <= '0';
      set_csum_begin_insert      <= '0';
      set_csum_rsvd_init         <= '0';
      set_txc_addr_0             <= '0';
      set_txc_addr_1             <= '0';
      set_txc_addr_2             <= '0';
      set_txc_addr_3             <= '0';
      set_txc_addr_4_n           <= '0';
      clr_txc_addr_3             <= '0';
      set_txcwr_rd_addr          <= '0';  --  sets the write side, read address to 0x0
      set_txcwr_wr_end           <= '0';  --  writes the end address to the memory in the next available location
      set_txc_en                 <= '0';  --  the enable bit to the write side of the memory
      set_txc_we                 <= '0';  --  the write enable bit to the write side of the memory
      inc_txd_addr_one           <= '0';
      set_txc_trdy               <= '0';
      init_bram                  <= '0';
      compare_addr2              <= '0';
      compare_addr0              <= '0';
      set_txc_trdy2              <= '0';
      clr_txc_trdy2              <= '0';
      enable_compare_addr0_cmplt <= '0';

      case txc_wr_cs is
        when TXC_ADDR2_WR =>
          set_txc_addr_2         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          txc_wr_ns              <= TXC_ADDR0_WR;
        when TXC_ADDR0_WR =>
          set_txc_addr_0         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          txc_wr_ns              <= WAIT_WR_CMPLT;
        when WAIT_WR_CMPLT =>
          set_txc_addr_0         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          set_txc_trdy2          <= '1';
          txc_wr_ns              <= TXC_WD0;
        when TXC_WD0 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' and
             (wrote_first_packet = '0' or txc_addr_3_dly = '1') then
            set_txc_addr_2         <= '1';  --Set the address to get the TxC Rd Address Pointer
            set_txc_en             <= '1';
            set_axi_flag           <= '1';
            clr_txc_addr_3         <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD1;
          else
            set_txc_addr_2         <= '0';  --Set the address to get the TxC Rd Address Pointer
            set_txc_en             <= '0';
            set_axi_flag           <= '0';
            clr_txc_addr_3         <= '0';
            compare_addr2          <= '0';
            txc_wr_ns              <= TXC_WD0;
          end if;

        when TXC_WD1 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_txc_trdy2          <= '0';
            set_csum_cntrl         <= '1';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD2;--WAIT_ADDR2_COMPARE_CMPLT;
          elsif axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '0' then
          -- need to force txc trdy HIGH since TVALID throttled
            set_txc_trdy2          <= '1';
            set_csum_cntrl         <= '0';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= WAIT_ADDR2_COMPARE_CMPLT;
          else
            set_txc_trdy2          <= '0';
            set_csum_cntrl         <= '0';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD1;
          end if;

        when WAIT_ADDR2_COMPARE_CMPLT =>
        -- now clear txc trdy to only allow a one clock pulse HIGH
          clr_txc_trdy2          <= '1';
          set_txc_addr_2         <= '1';
          set_txc_en             <= '1';
          compare_addr2          <= '1';
          txc_wr_ns              <= TXC_WD1;

        when TXC_WD2 =>
        -- Txc Tready has already been disabled
        --  wait for compare_addr2_cmplt, then
        --  set_txc_trdy2 will force axi_str_txc_tready_int_dly HIGH
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_csum_begin_insert      <= '1';
            set_txc_addr_2         <= '0';
            set_txc_en             <= '0';
            compare_addr2          <= '0';
            set_txc_trdy2          <= '0';
            txc_wr_ns                  <= TXC_WD3;
          else
            if axi_str_txc_tvalid_dly0 = '0'  or
               (txc_mem_full = '1' and axi_str_txc_tvalid_dly0 = '1') then
            --  If full wait for FULL and TVALID
            --  This will allow next elsif to be hit properly
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '1';
              set_txc_en             <= '1';
              compare_addr2          <= '1';
              set_txc_trdy2          <= '0';
              txc_wr_ns              <= TXC_WD2;


            elsif axi_str_txc_tvalid_dly0 = '1' and
              (compare_addr2_cmplt = '1' or compare_addr2_cmplt_dly = '1') then
              --  when full is '0', only need compare_addr2_cmplt to set set_txc_trdy2
              --    which will then allow this state to be exited to TXD_WD3
              --  when full is '1', then will need compare_addr2_cmplt_dly to to set set_txc_trdy2
              --    which will then allow this state to be exited to TXD_WD3
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '0';
              set_txc_en             <= '0';
              compare_addr2          <= '0';
              set_txc_trdy2          <= '1';
              txc_wr_ns                  <= TXC_WD2;
            else
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '1';
              set_txc_en             <= '1';
              compare_addr2          <= '1';
              set_txc_trdy2          <= '0';
              txc_wr_ns                  <= TXC_WD2;
            end if;
          end if;
        when TXC_WD3 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
          --  This is the earliest state to check for TxC FULL from TXC_WD0 state addr_2
          --  Register data, then assert full = 2 clks from rd
          --    Not FULL so write TxC Write Pointer to addr 0x3
            set_csum_rsvd_init         <= '1';
            txc_wr_ns                  <= TXC_WD4;
          else
            set_csum_rsvd_init         <= '0';
            txc_wr_ns                  <= TXC_WD3;
          end if;
        when TXC_WD4 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_txc_addr_0             <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            txc_wr_ns                  <= TXC_WD5;
          else
            set_txc_addr_0             <= '0';  --Set the address to get the TxD Rd Address Pointer
            set_txc_en                 <= '0';
            compare_addr0              <= '0';
            txc_wr_ns                  <= TXC_WD4;
          end if;
        when TXC_WD5 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' and axi_str_txc_tlast_dly0 = '1' then
            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '1';
            txc_wr_ns                  <= WAIT_ADDR0_COMPARE_CMPLT;
          else
            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '0';
            txc_wr_ns                  <= TXC_WD5;
          end if;
        when WAIT_ADDR0_COMPARE_CMPLT =>
          if compare_addr0_cmplt = '1' then
            set_txc_addr_1             <= '1'; -- this is one clock early, so do not set the we enable yet
            set_txc_en                 <= '1';
            set_txc_we                 <= '1';

            set_txc_addr_0             <= '0';
            set_txc_en                 <= '0';
            compare_addr0              <= '0';
            enable_compare_addr0_cmplt <= '0';
            txc_wr_ns                  <= WAIT_TXD_CMPLT;
          else
            set_txc_addr_1             <= '0';
            set_txc_en                 <= '0';
            set_txc_we                 <= '0';

            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '1';
            txc_wr_ns                  <= WAIT_ADDR0_COMPARE_CMPLT;
          end if;



        when WAIT_TXD_CMPLT =>
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1'  and
             axi_str_txd_tlast_dly0 = '1' then
            set_txc_addr_0        <= '0';
            set_txc_addr_1        <= '1';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WR_TXD_END_PNTR;
          elsif disable_txd_trdy_dly = '1' then
          -- Txd mem is full so get the current read pointer
          --  This can occure after tlast so check it in the following states
            set_txc_addr_0        <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_addr_1        <= '0';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_MEM;
          elsif update_bram_cnt(7) = '1'  then
          --Writing the current TxC write pointer so the read side can monitor it
            set_txc_addr_1        <= '1';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          else
            set_txc_addr_1        <= '0'; --Writing the current TxC write pointer so the read side can monitor it
            set_txc_addr_2        <= '0';
            set_txc_en            <= '0';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          end if;
        when WAIT_TXD_MEM =>
          if disable_txd_trdy_dly = '1' then
            -- Txd mem is full so get the current read pointer
            set_txc_addr_0        <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_addr_1        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_MEM;
          else
            set_txc_addr_0        <= '0';
            set_txc_addr_1        <= '1'; -- this is one clock early, so do not set the we enable yet
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          end if;
        when WR_TXD_END_PNTR =>
          if (load_data_1_dly = '1' and axi_str_txd_tlast_1 = '1' and tagmode_cross = "00") or 
          --  this condition is needed for packets less than 17 bytes and no tagging
            (axi_str_txd_tlast_1 = '1' and tagmode_cross /= "00" and tag_en_go = '0') then
            --  this condition is needed for packets less than 17 bytes and tagging
            inc_txd_addr_one      <= '0';
            set_txc_addr_4_n      <= '0'; -- Write the TxC End Value to address 0x4 - 0xn
            set_txc_en            <= '0';
            set_txc_we            <= '0';
            txc_wr_ns             <= WR_TXD_END_PNTR;
          else            
            inc_txd_addr_one      <= '1';
            set_txc_addr_4_n      <= '1'; -- Write the TxC End Value to address 0x4 - 0xn
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WR_TXC_PNTR;
          end if;
          
        when WR_TXC_PNTR =>
          if disable_txc_trdy_dly = '1' then
            set_txc_addr_0        <= '1';
            set_txc_addr_3        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';  
            set_txc_trdy          <= '0';
            txc_wr_ns             <= WR_TXC_PNTR;
          else          
            set_txc_addr_0        <= '0'; -- Write the TxC end pointer value to start the tx clint FSM
            set_txc_addr_3        <= '1';
            set_txc_en            <= '1';
            set_txc_we            <= '1';            
            set_txc_trdy          <= '1';
            txc_wr_ns             <= TXC_WD0;
          end if;          
          
--        when WR_TXC_PNTR =>
--            set_txc_addr_3        <= '1'; -- Write the TxC end pointer value to start the tx clint FSM
--            set_txc_addr_0        <= '0';
--            set_txc_en            <= '1';
--            set_txc_we            <= '1';
--            txc_wr_ns             <= TXC_WD0;
                    
        when others =>
          txc_wr_ns                <= TXC_ADDR2_WR;
      end case;
    end process;

    -----------------------------------------------------------------------------
    -- AXI Stream TX Control State Machine Sequencer
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXC_SEQ : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_wr_cs <= TXC_ADDR2_WR;
        else
          txc_wr_cs <= txc_wr_ns;
        end if;
      end if;
    end process;
    
    
    -----------------------------------------------------------------------------
    -- Needed to advance TxC FSM from write_txd_end_pntr state when tagmode_cross /= "00"
    -----------------------------------------------------------------------------
    TXC_GO_NO_TAG : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        tag_en_go <= set_tag_en_go;
      end if;
    end process;
        
    


    -----------------------------------------------------------------------------
    -- Delay the last write to TxC memory of the first packet after reset
    -----------------------------------------------------------------------------
    TX_INIT_INDICATOR_DLYS : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_addr_3_dly2 <= '0';
          txc_addr_3_dly3 <= '0';
        else
          txc_addr_3_dly2 <= txc_addr_3_dly;
          txc_addr_3_dly3 <= txc_addr_3_dly2;
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    -- Use above delay to hold off Tx Client FSM from starting until all
    --    TxD and TxC pointer information has been written to memory
    --
    --    This signal goes through a clock crossing circuit before it is
    --      registered in the Tx Client clock domain and used to start the
    --      Tx Client Read FSM
    -----------------------------------------------------------------------------
    TX_INIT_INDICATOR : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          tx_init_in_prog_int <= '1';
        else
          if txc_addr_3_dly3 = '1' then
            tx_init_in_prog_int <= '0';
          else
            tx_init_in_prog_int <= tx_init_in_prog_int;
          end if;
        end if;
      end if;
    end process;

    tx_init_in_prog <= tx_init_in_prog_int;

    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_1_TXD_WR_PNTR : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_1 = '1' then
          txc_addr_1 <= '1';
        else
          txc_addr_1 <= '0';
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_3_DELAY : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' or clr_txc_addr_3 = '1' then
          txc_addr_3_dly  <= '0';
        elsif set_txc_addr_3 = '1' then
          txc_addr_3_dly <= '1';
        else
          txc_addr_3_dly <= txc_addr_3_dly;
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    --  Generate address that will hold the End Address
    -----------------------------------------------------------------------------
    TXC_WR_ADDR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_mem_wr_addr      <= txc_min_wr_addr;
          txc_mem_wr_addr_last <= txc_wr_addr3;
          txc_mem_wr_addr_0    <= txc_wr_addr5;
          txc_mem_wr_addr_1    <= txc_wr_addr6;
        else
          if set_txc_addr_3 = '1' then
            --  increment the address for the next packet
            --  use the delayed signal to increment after the current address
            --  can be written
            if txc_mem_wr_addr = txc_max_wr_addr then
              --  if the max address is reached, loop to address 0x4
              txc_mem_wr_addr      <= txc_mem_wr_addr_0;
              txc_mem_wr_addr_last <= txc_wr_addr3;
              txc_mem_wr_addr_0    <= txc_mem_wr_addr_1;  --plus1
              txc_mem_wr_addr_1    <= txc_wr_addr6;       --plus2
            else
              --  otherwise just increment it
              txc_mem_wr_addr      <= txc_mem_wr_addr_0;
              txc_mem_wr_addr_last <= txc_mem_wr_addr;
              txc_mem_wr_addr_0    <= txc_mem_wr_addr_1;
              txc_mem_wr_addr_1    <= std_logic_vector(unsigned(txc_mem_wr_addr_1) + 1);
            end if;
          else -- Hold the current address until something changes
            txc_mem_wr_addr      <= txc_mem_wr_addr;
            txc_mem_wr_addr_last <= txc_mem_wr_addr_last;
            txc_mem_wr_addr_0    <= txc_mem_wr_addr_0;
            txc_mem_wr_addr_1    <= txc_mem_wr_addr_1;
          end if;
        end if;
      end if;
    end process;




    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_0_DELAY : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        txc_addr_0_dly1 <= set_txc_addr_0;
        txc_addr_0_dly2 <= txc_addr_0_dly1;
      end if;

    end process;


    -----------------------------------------------------------------------------
    --  Generate address that will hold the End Address
    -----------------------------------------------------------------------------
    MEM_TXC_WR_ADDR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then

        if set_txc_addr_4_n = '1' and set_txc_we = '1' then
          -- Provide the address for the End of packet address
          Axi_Str_TxC_2_Mem_Addr_int <= txc_mem_wr_addr;
        elsif set_txc_addr_3 = '1' and set_txc_we = '1' then
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr3; --set txc wr pointer
        elsif txc_addr_2 = '1' and  (txc_we = '0' or init_bram = '1') then
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr2; --get txc rd pointer
        elsif set_txc_addr_0 = '1' and (set_txc_we = '0' or init_bram = '1') then
          --  Monitor the read pointer for a full
          --  condition in the TxD Memory
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr0;
        elsif set_txc_addr_1 = '1' then
          --  Set the TxD write pointer to
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr1;
        else
          Axi_Str_TxC_2_Mem_Addr_int <= (others => '0');
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_Addr <= Axi_Str_TxC_2_Mem_Addr_int;
    txc_mem_wr_addr_plus1  <= txc_mem_wr_addr_0;
    txc_mem_wr_addr_plus2  <= txc_mem_wr_addr_1;

    -----------------------------------------------------------------------------
    --  This process remaps the strobe signal to the byte address offset minus
    --  one byte.
    -----------------------------------------------------------------------------
    END_ADDRESS_BYTE_OFFSET : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txD = '1' then
          end_addr_byte_offset <= (others => '0');
        elsif axi_str_txd_tlast_dly0 = '1' and axi_str_txd_tvalid_dly0 = '1' and 
              axi_str_txd_tready_int_dly = '1' then
          case axi_str_txd_tstrb_dly0 is
            when "1111" => end_addr_byte_offset <= "11";
            when "0111" => end_addr_byte_offset <= "10";
            when "0011" => end_addr_byte_offset <= "01";
            when others => end_addr_byte_offset <= "00";
          end case;
        else
          end_addr_byte_offset <= end_addr_byte_offset;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_WR_ADDR_VALUE : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' or init_bram = '1' then
          Axi_Str_TxC_2_Mem_Din_int <= (others => '0');
        elsif set_txc_addr_4_n = '1' then
        --write the ending address of the packet to memory minus one byte
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd_2 & axi_str_txd_2_mem_addr_int & end_addr_byte_offset;
        elsif set_txc_addr_3 = '1' then
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txc & txc_mem_wr_addr;
        else
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd & axi_str_txd_2_mem_addr_int_plus1;
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_Din <= Axi_Str_TxC_2_Mem_Din_int;

  --  Axi_Str_TxC_2_Mem_En  <= '1';
    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if (set_txc_en = '1' and set_txc_addr_2 = '0') or
           addr_2_en = '1' or init_bram = '1' then
          Axi_Str_TxC_2_Mem_En <= '1';
        else
          Axi_Str_TxC_2_Mem_En <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_WR_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_we = '1' then
          Axi_Str_TxC_2_Mem_We_int(0) <= '1';
        else
          Axi_Str_TxC_2_Mem_We_int(0) <= '0';
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_We <= Axi_Str_TxC_2_Mem_We_int;


    -----------------------------------------------------------------------------
    --  Delay set_txc_addr_2 to align with data
    -----------------------------------------------------------------------------
    TXC_ADDR2_DLY : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_2 = '1' then
          txc_addr_2  <= set_txc_addr_2;
        else
          txc_addr_2  <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay set_txc_we to align with address
    -----------------------------------------------------------------------------
    TXC_WE_DLY : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_we = '1' then
          txc_we  <= set_txc_we;
        else
          txc_we  <= '0';
        end if;
        txc_we_dly1 <= txc_we;
        txc_we_dly2 <= txc_we_dly1;

      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay set_txc_we to align with address
    -----------------------------------------------------------------------------
    ADDR2_MEM_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_2 = '1' and  set_txc_en = '1' then
          addr_2_en  <= set_txc_en;
        else
          addr_2_en  <= '0';
        end if;
        addr_2_en_dly1 <= addr_2_en;
        addr_2_en_dly2 <= addr_2_en_dly1;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Get the read pointer to check for FULL
    --  With ASYNC BRAM clock cannot read/write same address in memory at same
    --  time unless timing is met, so read until data matches
    -----------------------------------------------------------------------------
    MEM_TXC_RD_ADDR_PNTR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_rd_addr2_pntr_1 <= (others => '0');
          txc_rd_addr2_pntr   <= txc_min_wr_addr;
          compare_addr2_cmplt <= '0';
          compare_addr2_cmplt_dly <= '0';
        else

          if set_txc_addr_2 = '1' and addr_2_en_dly2 = '1' and txc_we_dly2 = '0' then
            txc_rd_addr2_pntr_1 <= Axi_Str_TxC_2_Mem_Dout(c_TxC_addrb_width -1 downto 0);

            if Axi_Str_TxC_2_Mem_Dout(c_TxC_addrb_width -1 downto 0) = txc_rd_addr2_pntr_1  and
               compare_addr2_cmplt = '0' then
              txc_rd_addr2_pntr   <= txc_rd_addr2_pntr_1;
              compare_addr2_cmplt <= '1';
            else
              txc_rd_addr2_pntr   <= txc_rd_addr2_pntr;
              compare_addr2_cmplt <= '0';
            end if;

          else
            txc_rd_addr2_pntr_1 <= txc_rd_addr2_pntr_1;
            txc_rd_addr2_pntr   <= txc_rd_addr2_pntr;
            compare_addr2_cmplt <= '0';
          end if;
          compare_addr2_cmplt_dly <= compare_addr2_cmplt;

        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Full flag indicator
    --    Does not begin comparison until 1st packet is written to memory
    -----------------------------------------------------------------------------
    TXC_FULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txc = '1' then
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
        elsif txc_mem_full = '1' and
           compare_addr2_cmplt = '1' and compare_addr2_cmplt_dly = '0' then
           --increments after it goes full, so use txc_mem_wr_addr for compare
          if txc_mem_wr_addr /= txc_rd_addr2_pntr then
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
          else
            txc_mem_full     <= txc_mem_full;
            txc_mem_not_full <= txc_mem_not_full;
          end if;
        elsif set_txc_addr_3 = '1' and set_txc_we = '1' then
          if txc_mem_wr_addr_plus1 = txc_rd_addr2_pntr then
            txc_mem_full     <= '1';
            txc_mem_not_full <= '0';
          else
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
          end if;
        else
          txc_mem_full     <= txc_mem_full;
          txc_mem_not_full <= txc_mem_not_full;
        end if;
      end if;
    end process;

    TXC_AFULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if txc_mem_wr_addr_plus2 = txc_rd_addr2_pntr then
          txc_mem_afull     <= '1';
        else
          txc_mem_afull     <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Throttle AXI Stream TxC
    --    Do not assert unless TxD is not in progress and the memory can
    --    accept data
    -----------------------------------------------------------------------------
    TXC_READY : process(AXI_STR_TXD_ACLK)
    begin



      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txc = '1' or clr_txc_trdy = '1' or clr_txc_trdy2 = '1' or
             set_txd_rdy = '1' or (txd_rdy = '1' and clr_txd_rdy = '0') or disable_txc_trdy = '1' or
             (AXI_STR_TXC_TLAST = '1' and AXI_STR_TXC_TVALID = '1' and axi_str_txc_tready_int = '1') or
             (compare_addr2 = '1' and axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1') then --do not need compare_addr0 because will clr at TLAST
          axi_str_txc_tready_int <= '0';
        else

          if txc_addr_3_dly = '1' then
            if (txc_mem_wr_addr = txc_rd_addr2_pntr and txc_mem_full = '1') then
              axi_str_txc_tready_int <= '0';
            elsif txc_mem_wr_addr = txc_rd_addr2_pntr and
                Axi_Str_TxC_2_Mem_We_int(0) = '1' then
              axi_str_txc_tready_int <= '0';
            else
              axi_str_txc_tready_int <= axi_str_txc_tready_int;
            end if;
          elsif set_txc_trdy = '1' then
            axi_str_txc_tready_int <= '1';
          elsif set_txc_trdy2 = '1' then
          --  need to force it high after address compare and after reset
            axi_str_txc_tready_int <= '1';
          else
            axi_str_txc_tready_int <= axi_str_txc_tready_int;
          end if;
        end if;
        axi_str_txc_tready_int_dly <= axi_str_txc_tready_int;
      end if;
    end process;

    AXI_STR_TXC_TREADY <= axi_str_txc_tready_int;  --fix me  need to look at all txc control and TDX tlast

    -----------------------------------------------------------------------------
    --  Register and hold the axi_flag information and CSUM Control information
    --    axi_flag
    --      0x5 = Status control
    --      0xA = Normal control
    --      0xF = Null Control
    --    CSUM
    --      00 = No CSUM will be performed
    --      01 = Partial Checksum will be performed
    --      10 = Full checksum offloading will be performed
    -----------------------------------------------------------------------------
    CNTRL_WD0 : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          axi_flag   <= (others => '0');
        elsif set_axi_flag = '1' then
          axi_flag   <= axi_str_txc_tdata_dly0(31 downto 28);
        else
          axi_flag   <= axi_flag;
        end if;
      end if;
    end process;

    enable_newFncEn <= '1' when axi_flag = "1010" else '0';

    CNTRL_WD1 : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          csum_cntrl <= (others => '0');
        elsif set_csum_cntrl = '1' then
          csum_cntrl <= axi_str_txc_tdata_dly0 (1 downto  0);
        else
          csum_cntrl <= csum_cntrl;
        end if;
      end if;
    end process;

      ---------------------------------------------------------------------------
      --  Delay signal to load csum value in csum calculation
      ---------------------------------------------------------------------------
      CHECK_FULL_SIG : process(AXI_STR_TXC_ACLK)
      begin

        if rising_edge(AXI_STR_TXC_ACLK) then
          check_full <= set_txc_addr_4_n;
        end if;
      end process;



    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Data Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXD_CONTROL : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_tvalid_dly0 <= '0';
          axi_str_txd_tlast_dly0  <= '0';
          clr_txd_trdy            <= '0';
        else
          axi_str_txd_tvalid_dly0 <= AXI_STR_TXD_TVALID;
          axi_str_txd_tlast_dly0  <= AXI_STR_TXD_TLAST;
          if axi_str_txd_tvalid = '1' and axi_str_txd_tlast = '1' and axi_str_txd_tready_int = '1' then
            clr_txd_trdy <= '1';
          else
            clr_txd_trdy <= '0';
          end if;
        end if;
      end if;
    end process;

    AXI_STR_TXD_TREADY <= axi_str_txd_tready_int;  --fix me  need to look at all txd control and TXC tlast

    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Data Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXD_IN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_tstrb_dly0  <= AXI_STR_TXD_TSTRB;
        axi_str_txd_tdata_dly0  <= AXI_STR_TXD_TDATA;
      end if;
    end process;


    DATA_REG_1 : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_all_hits = '1' then
          axi_str_txd_data_1  <= (others => '0');
          axi_str_txd_tstrb_1 <= (others => '0');
          axi_str_txd_tlast_1 <= '0';
        else
          if load_data_1 = '1' then
            axi_str_txd_data_1  <= axi_str_txd_tdata_dly0;
            axi_str_txd_tstrb_1 <= axi_str_txd_tstrb_dly0;
            axi_str_txd_tlast_1 <= axi_str_txd_tlast_dly0;
          else
            axi_str_txd_data_1  <= axi_str_txd_data_1;
            axi_str_txd_tstrb_1 <= axi_str_txd_tstrb_1;
            axi_str_txd_tlast_1 <= axi_str_txd_tlast_1;
          end if;
        end if;
      end if;
    end process;
    
    --  Needed for packets which are less than 17 bytes
    LOAD_TLAST_1_DLY : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        load_data_1_dly <= load_data_1;
      end if;
    end process;    

    DATA_REG_2 : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_all_hits = '1' then
          axi_str_txd_data_2  <= (others => '0');
          axi_str_txd_tstrb_2 <= (others => '0');
          axi_str_txd_tlast_2 <= '0';
        else
          if load_data_2 = '1' then
            axi_str_txd_data_2  <= axi_str_txd_tdata_dly0;
            axi_str_txd_tstrb_2 <= axi_str_txd_tstrb_dly0;
            axi_str_txd_tlast_2 <= axi_str_txd_tlast_dly0;
          else
            axi_str_txd_data_2  <= axi_str_txd_data_2;
            axi_str_txd_tstrb_2 <= axi_str_txd_tstrb_2;
            axi_str_txd_tlast_2 <= axi_str_txd_tlast_2;
          end if;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay the data one more clock for BRAM
    -----------------------------------------------------------------------------
    REG_TXD_DLY0 : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
          if set_mux_trans = '1' and set_mux_data_1_reg = '1' then
            axi_str_txd_tdata_dly1  <= transReg(7 downto 0) &
                                       axi_str_txd_data_1(23 downto 20) & transReg(11 downto 8) &
                                       axi_str_txd_data_1(15 downto  0);

          elsif set_mux_trans = '1' then
            axi_str_txd_tdata_dly1  <= transReg(7 downto 0) &
                                       axi_str_txd_tdata_dly0(23 downto 20) & transReg(11 downto 8) &
                                       axi_str_txd_tdata_dly0(15 downto  0);
          elsif set_mux_tag = '1' then
            axi_str_txd_tdata_dly1  <= newTagData_cross( 7 downto  0) & newTagData_cross(15 downto  8) &
                                       newTagData_cross(23 downto 16) & newTagData_cross(31 downto 24);
          elsif set_mux_data_1_reg = '1' then
            axi_str_txd_tdata_dly1  <= axi_str_txd_data_1;
          elsif set_mux_data_2_reg = '1' then
            axi_str_txd_tdata_dly1  <= axi_str_txd_data_2;
          elsif set_mux_dly = '1' then
            axi_str_txd_tdata_dly1  <= axi_str_txd_tdata_dly0;
          elsif axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
            axi_str_txd_tdata_dly1  <= axi_str_txd_tdata_dly0;
          else
            axi_str_txd_tdata_dly1  <= axi_str_txd_tdata_dly1;
          end if;
      end if;
    end process;

    vlan_sel <= tag0TotalHit & newTagTotalHit & transTotalHit;

    -----------------------------------------------------------------------------
    --  AXI Stream TX Data State Machine - combinational/combinatorial
    --    Used to provide the control to write the data to the BRAM
    --    This state machine will throttle the Transmit AXI Stream Control state
    --      machine until after the data information has been received.
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXD_CMB : process (txd_wr_cs,axi_str_txd_tvalid_dly0,
      axi_str_txd_tlast_dly0,
      axi_str_txd_tstrb_dly0,wrote_first_packet,axi_str_txd_tready_int_dly,
      txd_rd_pntr,txd_mem_full,txd_mem_afull,update_cnt,
      txd_rd_pntr_hold,free_up_memory,txd_max_wr_addr_minus10,txd_mem_clr_words,
      decode_dly4,vlan_sel,axi_str_txd_tstrb_1,txd_rd_pntr_hold_plus3,txd_rd_pntr_hold_plus9,
      axi_str_txd_tstrb_2,axi_str_txd_tlast_1,axi_str_txd_tlast_2,
      txd_throttle_dly,ignore_tvalid_dly,compare_addr0_cmplt,ignore_txd_tvalid,
      axi_str_txd_2_mem_addr_int,txd_max_wr_addr,nine,
      check_full,txd_max_wr_addr_minus4,tagmode_cross)
    begin

      inc_txd_wr_addr     <= '0';
      set_txd_we          <= "0000";
      set_txd_en          <= '0';
      set_first_packet    <= '0';
      set_txd_rdy         <= '0';
      clr_txd_rdy         <= '0';
      clr_full_pntr       <= '0';
      disable_txd_trdy    <= '0';
      disable_txc_trdy    <= '0';
      halt_pntr_update    <= '0';
      set_mux_dly         <= '0';
      clr_mux_dly         <= '0';
      set_vlan_bram_en    <= '0';
      clr_vlan_bram_en    <= '0';
      txd_throttle        <= '0';
      clr_all_hits        <= '0';
      set_txd_tlast_rcvd  <= '0';
      setCheckTag0Tpid    <= '0';
      setCheckTag1Tpid    <= '0';
      set_mux_tag         <= '0';
      set_mux_trans       <= '0';
      set_mux_data_1_reg  <= '0';
      set_mux_data_2_reg  <= '0';
      ignore_txd_trdy     <= '0';
      load_data_1         <= '0';
      load_data_2         <= '0';
      ignore_tvalid       <= '0';
      set_ignore_txd_tvalid <= '0';

      update_rd_pntrs     <= '0';
      set_decode_dly      <= '0';
      
      inhibit_checktag0tpid <= '0';
      set_tag_en_go       <= '0';





      case txd_wr_cs is
        when IDLE =>
          if compare_addr0_cmplt = '1' then
          --  Requirement is that the TXD and TXC interfaces use the same clock
          --    so it is OK to used the TXC signals in the TXD state machine
            set_txd_rdy <= '1';
            txd_wr_ns   <= TXD_PRM;
          else
            set_txd_rdy <= '0';
            txd_wr_ns   <= IDLE;
          end if;

        when TXD_PRM =>
--      Made change to ensure TxD Memory is never full here.
--      The memory can always accept data at the start of a transfer
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
          --  delay incrementing pointer until next data
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            set_mux_dly         <= '1';
            txd_wr_ns           <= DST_SRC;
          else
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_mux_dly         <= '0';
            txd_wr_ns           <= TXD_PRM;
          end if;

        when DST_SRC =>
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
            inc_txd_wr_addr     <= '1';
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            clr_mux_dly         <= '1';
            set_vlan_bram_en    <= '0';
            txd_throttle        <= '0';
            txd_wr_ns           <= SRC;
          else
            inc_txd_wr_addr     <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            clr_mux_dly         <= '0';
            set_vlan_bram_en    <= '0';
            txd_throttle        <= '0';
            txd_wr_ns           <= DST_SRC;
          end if;
        when SRC =>
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
            -- no vlan
            --  can never have a case of all zeroes here since this is the T/L field
            inc_txd_wr_addr     <= '1';
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            clr_txd_rdy         <= '0';
            disable_txd_trdy    <= '0';

            set_vlan_bram_en    <= '1'; 
            clr_vlan_bram_en    <= '0'; 
            txd_throttle        <= '1';
            setCheckTag0Tpid    <= '1'; 
            txd_wr_ns           <= VLAN1;
          else
            inc_txd_wr_addr     <= '0';
            set_vlan_bram_en    <= '0';
            txd_throttle        <= '0';
            txd_wr_ns           <= SRC;
          end if;
        when VLAN1 =>
          if (axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1') or
          ignore_tvalid_dly = '1' then
          --do not increment address and exit this state until axi_str_txd_tready_int_dly = '1'
            clr_vlan_bram_en    <= '0';
            inc_txd_wr_addr     <= '1';

            txd_throttle        <= '1';
            setCheckTag1Tpid    <= '1';
            ignore_txd_trdy     <= '1';
            load_data_1         <= '1';
            set_vlan_bram_en    <= '1';
            txd_wr_ns           <= VLAN2;
          else
          -- axi_str_txd_tvalid_dly0 = '0' so wait for valid data
            inhibit_checktag0tpid <= '1';
            clr_vlan_bram_en    <= '0';
            inc_txd_wr_addr     <= '0';
            txd_throttle        <= '1';
            setCheckTag1Tpid    <= '0';
            ignore_txd_trdy     <= '1';
            load_data_1         <= '0';
            set_vlan_bram_en    <= '0';  -- 0510_2011
            txd_wr_ns           <= WAIT_TVALID;
          end if;

        when WAIT_TVALID =>
          if txd_throttle_dly = '0' then
          --Return the VLAN1 1 clock after txd_throttle is asserted LOW
          --this ensures axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1'
          --so FSM will not return back to this state
            clr_vlan_bram_en    <= '0';
            inc_txd_wr_addr     <= '0';

            txd_throttle        <= '1';
            setCheckTag0Tpid    <= '1';
            setCheckTag1Tpid    <= '0';
            ignore_txd_trdy     <= '1';
            load_data_1         <= '0';
            set_vlan_bram_en    <= '1';
            ignore_tvalid       <= '1';
            txd_wr_ns           <= VLAN1;
          elsif axi_str_txd_tvalid_dly0 = '1' then
          --Wait for tvalid to assert, then pulse throttle low for 1 clock cycle
            clr_vlan_bram_en    <= '0';
            inc_txd_wr_addr     <= '0';

            txd_throttle        <= '0';
            setCheckTag0Tpid    <= '1';
            setCheckTag1Tpid    <= '0';
            ignore_txd_trdy     <= '1';
            load_data_1         <= '0';
            set_vlan_bram_en    <= '1';
            ignore_tvalid       <= '0';
            txd_wr_ns           <= WAIT_TVALID;
          else
            clr_vlan_bram_en    <= '0';
            inc_txd_wr_addr     <= '0';

            txd_throttle        <= '1';
            setCheckTag0Tpid    <= '0';
            setCheckTag1Tpid    <= '0';
            ignore_txd_trdy     <= '1';
            load_data_1         <= '0';
            set_vlan_bram_en    <= '0';  -- 0510_2011
            ignore_tvalid       <= '0';
            txd_wr_ns           <= WAIT_TVALID;
          end if;

        when VLAN2 =>
          if axi_str_txd_tlast_1 = '1' and tagmode_cross = "00" then --or           --  received TLAST (0-2 bytes) or
--             axi_str_txd_tstrb_1 /= "1111" then     --  all strobes were not set (end of packet)
          --  Received TLAST and this cannot be a VLAN TAG Frame,
          --  But it can TAG so see if tagmode_cross = "00".  
          --  If tagmode_cross ="00" then write data and wait for next packet.
          --  If tagmode_cross /="00" then do not write, must tag, then write data. 
            inc_txd_wr_addr     <= '0';
            disable_txd_trdy    <= '0';
            set_mux_data_1_reg  <= '1';
            set_txd_we          <= axi_str_txd_tstrb_1;
            set_txd_en          <= '1';
            txd_throttle        <= '1';
            clr_txd_rdy         <= '1';
            txd_wr_ns             <= WAIT_WR1;
          elsif axi_str_txd_tlast_1 = '1' and tagmode_cross /= "00" then 
          -- 0520_2011 added this condition
          --  Received TLAST and this cannot be a VLAN TAG Frame,
          --  But it can TAG a non VLAN frame so see if tagmode_cross = "00".  
          --  If tagmode_cross ="00" then write data and wait for next packet.
          --  If tagmode_cross /="00" then do not write, must tag, then write data. 
            inc_txd_wr_addr     <= '0';
            disable_txd_trdy    <= '0';
            set_mux_data_1_reg  <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            txd_throttle        <= '1';
            clr_txd_rdy         <= '1';
            set_decode_dly      <= '1';
            set_ignore_txd_tvalid <= '1';
            txd_wr_ns             <= DECODE;          
          elsif axi_str_txd_tvalid_dly0 = '1' then
            set_vlan_bram_en    <= '1';
            setCheckTag1Tpid    <= '1';
            set_decode_dly      <= '1';
            txd_throttle        <= '1';
            ignore_txd_trdy     <= '1';
            load_data_2         <= '1';
--            clr_vlan_bram_en    <= '1'; --mw 0510_2011
            txd_wr_ns           <= DECODE;
          else
-- 0510_2011 Moved below signals to above elseif.  Must be checked only when TVLAID is asserted          
-- 0510_2011          --   axi_str_txd_tvalid_dly0 = '0' so need to wait for valid data
-- 0510_2011          --  but set bram whil it is invalid so once it is valid it will be ready
-- 0510_2011            --100817
-- 0510_2011            set_vlan_bram_en    <= '1';
-- 0510_2011            setCheckTag1Tpid    <= '1';
            --100817

            set_vlan_bram_en    <= '0';            
            setCheckTag1Tpid    <= '0';            
            txd_throttle        <= '1';
            ignore_txd_trdy     <= '1';
            load_data_2         <= '0';
            clr_vlan_bram_en    <= '0';
            txd_wr_ns           <= VLAN2;
          end if;
        when DECODE =>
          if (axi_str_txd_tlast_2 = '1') then -- or --ignore tvalid
--              axi_str_txd_tstrb_2 /= "1111") then --ignore tvalid
            set_ignore_txd_tvalid <= '1';
          else
            set_ignore_txd_tvalid <= '0';
          end if;


          if (axi_str_txd_tvalid_dly0 = '1' and
              --  tlast did not occur in previous state and neither did
              axi_str_txd_tlast_2 = '0' and axi_str_txd_tstrb_2 = "1111") or

             (axi_str_txd_tlast_2 = '1' or
              axi_str_txd_tlast_1 = '1') then 
             
            if decode_dly4 = '1' then
              case vlan_sel is
                when "111" | "110" =>
                  txd_throttle        <= '0';
                  set_mux_tag         <= '1';
                  set_txd_we          <= "1111";
                  set_txd_en          <= '1';
                when "101" =>
                  txd_throttle        <= '0';
                  set_mux_trans       <= '0';
                  set_txd_we          <= "0000";
                  set_txd_en          <= '0';
                when "100"  =>
                  txd_throttle        <= '0';
                  set_mux_tag         <= '0';
                  set_txd_we          <= "0000";
                  set_txd_en          <= '0';
                when "010" | "011" =>
                  txd_throttle        <= '1';
                  set_mux_tag         <= '1';
                  set_txd_we          <= "1111";
                  set_txd_en          <= '1';
                when "001"  =>
                  txd_throttle        <= '0';
                  set_mux_trans       <= '1';
                  set_mux_data_1_reg  <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_1;
                  set_txd_en          <= '1';
                when others => --"000"
                  if axi_str_txd_tlast_1 = '1' then
                    txd_throttle        <= '0';
                    set_mux_data_1_reg  <= '1';
                    set_txd_we          <= axi_str_txd_tstrb_1;
                    set_txd_en          <= '1';
                  else
                    txd_throttle        <= '0';
                    set_mux_data_1_reg  <= '0';
                    set_txd_we          <= "0000";
                    set_txd_en          <= '0';
                  end if;
              end case;
              txd_wr_ns           <= STTR;
            else
              set_txd_we          <= "0000";
              set_txd_en          <= '0';
              set_mux_dly         <= '0';
              txd_throttle        <= '1';
              txd_wr_ns           <= DECODE;
            end if;
          else
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_mux_dly         <= '0';
            txd_throttle        <= '1';
            txd_wr_ns           <= DECODE;
          end if;
          ignore_txd_trdy     <= '1';
        when STTR =>
          if axi_str_txd_tvalid_dly0 = '1' or ignore_txd_tvalid = '1' then

            case vlan_sel is
              when "111" =>
                inc_txd_wr_addr     <= '1';
                set_mux_trans       <= '1';
                set_txd_we          <= axi_str_txd_tstrb_2;
                set_txd_en          <= '1';
                txd_throttle        <= '0';
                txd_wr_ns           <= TRANSLATE;
              when "110" =>
                inc_txd_wr_addr     <= '1';
                set_mux_data_2_reg  <= '1';
                set_txd_we          <= axi_str_txd_tstrb_2;
                set_txd_en          <= '1';
                txd_throttle        <= '0';
                txd_wr_ns           <= TAG;
              when "101"  =>  --**
                inc_txd_wr_addr     <= '0';
                set_mux_trans       <= '1';
                set_txd_we          <= "1111";
                set_txd_en          <= '1';
                txd_throttle        <= '0';
                txd_wr_ns           <= TRANSLATE;
              when "100"  =>
                inc_txd_wr_addr     <= '0';
                set_mux_data_2_reg  <= '0';
                set_txd_we          <= "0000";
                set_txd_en          <= '0';
                txd_throttle        <= '0';
                txd_wr_ns           <= STRIP;
              when "011"  =>
                inc_txd_wr_addr     <= '1';
                set_mux_data_1_reg  <= '1';
                set_mux_trans       <= '1';
                set_txd_we          <= axi_str_txd_tstrb_1;
                set_txd_en          <= '1';
                txd_throttle        <= '0';
                txd_wr_ns           <= TRANSLATE;
              when "010" =>
                inc_txd_wr_addr     <= '1';
                set_mux_data_1_reg  <= '1';
                set_txd_we          <= axi_str_txd_tstrb_1; --  first vlan strobes;
                set_txd_en          <= '1';
                txd_throttle        <= '0';
                txd_wr_ns           <= TAG;
              when "001" =>
                inc_txd_wr_addr     <= '1';
                set_mux_data_2_reg  <= '0';
                set_txd_we          <= "0000";
                set_txd_en          <= '0';
                txd_throttle        <= '0';
                txd_wr_ns           <= TRANSLATE;
              when others => --"000"
                if axi_str_txd_tlast_1 = '1' then
                -- added 0520_2011 - VALN_sel = "000" and axi_str_txd_tlast_1 = '1'
                --data was written in previous state, so exit
                  inc_txd_wr_addr     <= '0';
                  set_mux_data_1_reg  <= '0';
                  set_txd_we          <= "0000";
                  set_txd_en          <= '0';
                  txd_throttle        <= '0';
                  set_tag_en_go       <= '1';
                  txd_wr_ns           <= WAIT_WR1;                
                else
                  inc_txd_wr_addr     <= '0';
                  set_mux_data_1_reg  <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_1;
                  set_txd_en          <= '1';
                  txd_throttle        <= '0';
                  txd_wr_ns           <= TRANSLATE;
                end if;
            end case;
          else
            inc_txd_wr_addr     <= '0';
            set_mux_data_2_reg  <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            txd_throttle        <= '0';
            txd_wr_ns           <= STTR;
          end if;
          ignore_txd_trdy     <= '1';
        when STRIP =>
          if axi_str_txd_tvalid_dly0 = '1' or ignore_txd_tvalid = '1' then
            if axi_str_txd_tlast_2 = '1' then
              inc_txd_wr_addr     <= '0';
              set_mux_dly         <= '0';
              set_txd_we          <= axi_str_txd_tstrb_2; --  second vlan strobes
              set_txd_en          <= '1';
              clr_txd_rdy         <= '1';
              txd_wr_ns           <= WAIT_WR1;
            elsif axi_str_txd_tlast_dly0 = '1' then
              inc_txd_wr_addr     <= '0';
              set_mux_dly         <= '0';
              set_txd_we          <= axi_str_txd_tstrb_dly0;
              set_txd_en          <= '1';
              clr_txd_rdy         <= '1';
              txd_wr_ns           <= WAIT_WR1;
            else
              inc_txd_wr_addr     <= '0';
              set_mux_dly         <= '1';
              set_txd_we          <= axi_str_txd_tstrb_dly0;
              set_txd_en          <= '1';
              txd_wr_ns           <= TXD_WRT;
            end if;
          else
            inc_txd_wr_addr     <= '0';
            set_mux_dly         <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            txd_wr_ns           <= STRIP;
          end if;
        when TAG =>
          if axi_str_txd_tvalid_dly0 = '1' or ignore_txd_tvalid = '1' then
            case vlan_sel is
              when "010" =>
                if axi_str_txd_tlast_1 = '1' then
                  inc_txd_wr_addr     <= '0';
                  set_mux_data_2_reg  <= '0';
                  set_mux_dly         <= '0';
                  set_txd_we          <= "0000"; --  first vlan strobes
                  set_txd_en          <= '0';
                  clr_txd_rdy         <= '1';
                  set_tag_en_go       <= '1';  --added 0520_2011
                  txd_wr_ns           <= WAIT_WR1;
                elsif axi_str_txd_tlast_2 = '1' then --and axi_str_txd_tstrb_2 /= "0000" then
                  inc_txd_wr_addr     <= '1';
                  set_mux_data_2_reg  <= '1';
                  set_mux_dly         <= '0';
                  set_txd_we          <= axi_str_txd_tstrb_2; --  second vlan strobes
                  set_txd_en          <= '1';
                  txd_wr_ns           <= WAIT_STATE;
--                elsif axi_str_txd_tlast_2 = '1' or axi_str_txd_tstrb_2 = "0000" then
--                  inc_txd_wr_addr     <= '0';
--                  set_mux_data_2_reg  <= '0';
--                  set_mux_dly         <= '0';
--                  set_txd_we          <= "0000"; --  second vlan strobes
--                  set_txd_en          <= '0';
--                  clr_txd_rdy         <= '1';
--                  txd_wr_ns           <= WAIT_WR1;
                else
                  inc_txd_wr_addr     <= '1';
                  set_mux_data_2_reg  <= '0';
                  set_mux_dly         <= '1';
                  set_txd_we          <= "0000";
                  set_txd_en          <= '0';
                  txd_wr_ns           <= WAIT_STATE;
                end if;
              when others  => -- "110"
                if axi_str_txd_tlast_dly0 = '1' then
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '0';
                  set_txd_we          <= "0000"; --already wrote it --axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '0';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
                else
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '1';
                  set_txd_we          <= "0000";
                  set_txd_en          <= '0';
                  txd_wr_ns           <= TXD_WRT;
                end if;
            end case;
          else
            inc_txd_wr_addr     <= '0';
            set_mux_dly         <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            txd_wr_ns           <= TAG;
          end if;
        when TRANSLATE =>
          if axi_str_txd_tvalid_dly0 = '1' or ignore_txd_tvalid = '1' then
            case vlan_sel is
              when "111" =>  --**
                inc_txd_wr_addr     <= '1';
                set_mux_dly         <= '0';
                set_txd_we          <= "0000";
                set_txd_en          <= '0';
                txd_wr_ns           <= WAIT_STATE;
              when "101"  =>
                if axi_str_txd_tlast_dly0 = '1' then
                  inc_txd_wr_addr     <= '1';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
                else
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '1';
                  set_txd_we          <= "0000";
                  set_txd_en          <= '0';
                  txd_wr_ns           <= TXD_WRT;
                end if;
              when "011"  =>
                if axi_str_txd_tlast_2 = '1' then
                --CANNOT HAVE ALL ZERO STROBES HERE
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '0';
                  set_txd_we          <= "0000";
                  set_txd_en          <= '0';
                  txd_wr_ns           <= WAIT_STATE;
                else
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '1';
                  set_txd_we          <= "0000";
                  set_txd_en          <= '0';
                  txd_wr_ns           <= TXD_WRT;
                end if;
              when "001" =>
                set_mux_dly         <= '1';
                if axi_str_txd_tlast_dly0 = '1' or axi_str_txd_tlast_2 = '1' then
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
                else -- TLAST has not been received and neither have strobes of zeroes
                  inc_txd_wr_addr     <= '0';
                  set_txd_we          <= "1111";
                  set_txd_en          <= '1';
                  txd_wr_ns           <= TXD_WRT;
                end if;
              when others => --when "000" =>
                if axi_str_txd_tlast_2 = '1' then
                  inc_txd_wr_addr     <= '1';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
--                elsif axi_str_txd_tstrb_2 = "0000" then
--                  inc_txd_wr_addr     <= '0';
--                  set_mux_dly         <= '0';
--                  set_txd_we          <= axi_str_txd_tstrb_2;
--                  set_txd_en          <= '0';
--                  txd_wr_ns           <= WAIT_WR1;
                else
                  inc_txd_wr_addr     <= '1';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  txd_wr_ns           <= TXD_WRT;
                end if;
            end case;
          else
            inc_txd_wr_addr     <= '0';
            set_mux_dly         <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            txd_wr_ns           <= TRANSLATE;
          end if;
        when WAIT_STATE =>
          --Should only get to this state when vlan_sel = "010" ,"011", or "111"
          if axi_str_txd_tvalid_dly0 = '1' or ignore_txd_tvalid = '1' then
            case vlan_sel is
              when "010" =>
                if axi_str_txd_tlast_2 = '1' then
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '0';
                  set_txd_we          <= "0000";
                  set_txd_en          <= '0';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
                elsif axi_str_txd_tlast_dly0 = '1' then
                  inc_txd_wr_addr     <= '1';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
                else
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  txd_wr_ns           <= TXD_WRT;
                end if;
              when "011" => -- "011"
                if axi_str_txd_tlast_2 = '1' then
                  inc_txd_wr_addr     <= '1';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_2;
                  set_txd_en          <= '1';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
                elsif axi_str_txd_tlast_dly0 = '1' then
                  inc_txd_wr_addr     <= '1';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
                else
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  txd_wr_ns           <= TXD_WRT;
                end if;
              when others => -- "111"
                if axi_str_txd_tlast_2 = '1' then
                  inc_txd_wr_addr     <= '1';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_2;
                  set_txd_en          <= '1';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
                elsif axi_str_txd_tlast_dly0 = '1' then
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  clr_txd_rdy         <= '1';
                  txd_wr_ns           <= WAIT_WR1;
                else
                  inc_txd_wr_addr     <= '0';
                  set_mux_dly         <= '1';
                  set_txd_we          <= axi_str_txd_tstrb_dly0;
                  set_txd_en          <= '1';
                  txd_wr_ns           <= TXD_WRT;
                end if;
            end case;
          else
            inc_txd_wr_addr     <= '0';
            set_mux_dly         <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            txd_wr_ns           <= WAIT_STATE;
          end if;
        when  TXD_WRT =>
          if txd_mem_full = '1' and axi_str_txd_tready_int_dly = '0' then
          --memory is full when axi_str_txd_tready_int_dly = '0'
            inc_txd_wr_addr     <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_first_packet    <= '0';
            clr_txd_rdy         <= '0';
            disable_txd_trdy    <= '1';
            txd_wr_ns           <= MEM_FULL;
          elsif axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
            inc_txd_wr_addr     <= '1';
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            if axi_str_txd_tlast_dly0 = '1' then
              if wrote_first_packet = '0' then
                set_first_packet <= '1';
              else
                set_first_packet <= '0';
              end if;

              clr_txd_rdy         <= '1';
              disable_txc_trdy    <= '1';
              disable_txd_trdy    <= '0';
              clr_txd_rdy         <= '1';
              txd_wr_ns           <= WAIT_WR1;
            else
            --  received data (normal receive), so continue receiving data
              set_first_packet    <= '0';
              clr_txd_rdy         <= '0';
              disable_txd_trdy    <= '0';
              txd_wr_ns           <= TXD_WRT;
            end if;
          else
            inc_txd_wr_addr     <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_first_packet    <= '0';
            clr_txd_rdy         <= '0';
            disable_txd_trdy    <= '0';
            txd_wr_ns           <= TXD_WRT;
          end if;
       when MEM_FULL =>
          --  stay here until the read pointer updates by 4 words or more.  The read side operates on bytes,
          --  the write side operates on words.
          --    The read pointer updates every 512 bytes (128 words) and at the end of a packet.
          --      The samallest packet the can be sent is 15bytes, but since the BRAM is 32 bit aligned,
          --      the read side will usually update the read pointer by a minimum of 16 bytes (4 words).  However,
          --      it can update by by less than 16 bytes (4 words).  This can occure if a packet started at read
          --      address 0x1A4 (write address 0x69), and the packet is 516 bytes in length (129 words).  Here the read pointer
          --      will update at 0x3A4 (write address 0xE9 - 128 words) then again at the end of the packet at 0x3A8
          --      (write address 0xEA).
          --        If this occures the below logic will detect it and update the read pointer, but stay in this
          --        state until the next update occurs.  The next update is guaranteed to be greater than 4 words,
          --        which will allow the full pointers to be cleared for the next packet.
          inc_txd_wr_addr     <= '0';
          set_txd_we          <= "0000";
          set_txd_en          <= '0';
          set_first_packet    <= '0';
          clr_txd_rdy         <= '0';
          if txd_rd_pntr = txd_rd_pntr_hold then
          --  stay here until an update occurs
            update_rd_pntrs  <= '0';
            disable_txd_trdy <= '1';
            clr_full_pntr    <= '0';
            txd_wr_ns        <= MEM_FULL;
          else
          --  The read pointer was updated to determine if it was updated by 4 words or more
          --    If not, update the hold pointers, but stay in this state
            if txd_rd_pntr_hold <= txd_max_wr_addr_minus4 then
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x0 - 0x1FB
              if txd_rd_pntr > txd_rd_pntr_hold_plus3 then
              -- an update of 4 words or greater occured so exit this state
                update_rd_pntrs  <= '0';
                disable_txd_trdy <= '0';
                clr_full_pntr    <= '1';
                txd_wr_ns        <= TXD_WRT;
              else
              --  the update was less than 4 words
              --    (txd_rd_pntr <= txd_rd_pntr_hold_plus3)
                if txd_rd_pntr < txd_rd_pntr_hold then
                --  the read pointer wrapped, so exit because the update was > 4 words
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              end if;
            else
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x1FC- 0x1FF
              if txd_rd_pntr_hold_plus3 = txd_max_wr_addr then
              --  txd_rd_pntr = 0x1FC for 2048 byte memory, so txd_rd_pntr_hold_plus3 = max memory size
                if (txd_rd_pntr <= txd_rd_pntr_hold) then
                --  the update was >= 4 words so exit
                --    for a 2048 memory, txd_rd_pntr_hold = 0x1FC
                --      if txd_rd_pntr is between 0x0 and 0x1FB then an update of 4 or more words occurred
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              else
              --  txd_rd_pntr = 0x1FD, 0x1FE, or 0x1FF for 2048 byte memory,
              --  so the minimum txd_rd_pntr_hold_plus3 can be is 0, 1, or 2
                if (txd_rd_pntr > txd_rd_pntr_hold_plus3) and (txd_rd_pntr < txd_rd_pntr_hold) then
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr has to be tween 0x1 and 0x1FC to exit this state
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr has to be tween 0x2 and 0x1FD to exit this state
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr has to be tween 0x3 and 0x1FE to exit this state
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  txd_rd_pntr did not update by 4 or more words, so update hold poointers and stay in this state
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited BUT
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr was only updated 1-3 words to 0x1FE, 0x1FF, or 0x0, so stay here
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr was only updated 1-3 words to 0x1FF, 0x0, or 0x1, so stay here
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr was only updated 1-3 words to 0x0, 0x1, or 0x2, so stay here
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              end if;
            end if;
          end if;

        when WAIT_WR1 =>
          disable_txc_trdy  <= '1';
          disable_txd_trdy  <= '0';

          if check_full = '1' then
            txd_wr_ns         <= WAIT_WR2;
          else
            txd_wr_ns         <= WAIT_WR1;
          end if;
        when WAIT_WR2 =>
          if txd_mem_clr_words = '1' then
            disable_txc_trdy  <= '1';
            disable_txd_trdy  <= '1';
            txd_wr_ns         <= CLR_WORDS;
          else
            if wrote_first_packet = '0' then
              set_first_packet <= '1';
            else
              set_first_packet <= '0';
            end if;
            clr_all_hits      <= '1';
            clr_txd_rdy       <= '0';

            disable_txc_trdy  <= '0';
            disable_txd_trdy  <= '0';
            txd_wr_ns         <= IDLE;
          end if;
        when CLR_WORDS =>
          --  stay here until the read pointer updates by 10 words or more.  The read side operates on bytes,
          --  the write side operates on words.
          --    The read pointer updates every 512 bytes (128 words) and at the end of a packet.
          --      The samallest packet the can be sent is 15bytes, but since the BRAM is 32 bit aligned,
          --      the read side will usually update the read pointer by a minimum of 16 bytes (4 words).  However,
          --      it can update by by less than 16 bytes (4 words).  This can occure if a packet started at read
          --      address 0x1A4 (write address 0x69), and the packet is 516 bytes in length (129 words).  Here the read pointer
          --      will update at 0x3A4 (write address 0xE9 - 128 words) then again at the end of the packet at 0x3A8
          --      (write address 0xEA).
          --        If this occures the below logic will detect it and update the read pointer, but stay in this
          --        state until the next update occurs.  The next update is guaranteed to be greater than 10 words,
          --        which will allow the full pointers to be cleared for the next packet.
          inc_txd_wr_addr     <= '0';
          set_txd_we          <= "0000";
          set_txd_en          <= '0';
          set_first_packet    <= '0';
          clr_txd_rdy         <= '0';

          if update_cnt <= nine then
            if txd_rd_pntr = txd_rd_pntr_hold then
            --  stay here until an update occurs
              update_rd_pntrs  <= '0';
              halt_pntr_update <= '1';
              disable_txc_trdy <= '1';
              disable_txd_trdy <= '1';
              clr_full_pntr    <= '0';
              txd_wr_ns        <= CLR_WORDS;
            else
            --  The read pointer was updated to determine if it was updated by 10 words or more
            --    If not, update the hold pointers, but stay in this state
              if txd_rd_pntr_hold <= txd_max_wr_addr_minus10 then
              --  for 2048 mem this covers from txd_rd_pntr_hold = 0x0 - 0x1F5
                if txd_rd_pntr > txd_rd_pntr_hold_plus9 then
                -- an update of 10 words or greater occured so exit this state
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_all_hits     <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  the update was less than 10 words
                --    (txd_rd_pntr <= txd_rd_pntr_hold_plus9)
                  if txd_rd_pntr < txd_rd_pntr_hold then
                  --  the read pointer wrapped, so exit because the update was > 10 words
                    if wrote_first_packet = '0' then
                      set_first_packet <= '1';
                    else
                    --  the update was less than 10 words, so update the read hold pointers and stay here until the next update
                    --    txd_rd_pntr >= txd_rd_pntr_hold
                      set_first_packet <= '0';
                    end if;
                    update_rd_pntrs  <= '0';
                    halt_pntr_update <= '0';
                    disable_txd_trdy <= '0';
                    clr_full_pntr    <= '1';
                    clr_all_hits     <= '1';
                    clr_txd_rdy      <= '0';
                    txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                  else
                  --  the update was less than 10 words, so update the read hold pointers and stay here until the next update
                  --    txd_rd_pntr >= txd_rd_pntr_hold
                    update_rd_pntrs  <= '1';
                    halt_pntr_update <= '1';
                    disable_txc_trdy <= '1';
                    disable_txd_trdy <= '1';
                    clr_full_pntr    <= '0';
                    txd_wr_ns        <= CLR_WORDS;
                  end if;
                end if;

              else
                --  for 2048 mem this covers from txd_rd_pntr_hold = 0x1F6- 0x1FF
                if txd_rd_pntr_hold_plus9 = txd_max_wr_addr then
                --  txd_rd_pntr = 0x1F6 for 2048 byte memory, so txd_rd_pntr_hold_plus9 = max memory size
                  if (txd_rd_pntr <= txd_rd_pntr_hold) then
                  --  the update was >= 10 words so exit
                  --    for a 2048 memory, txd_rd_pntr_hold = 0x1F6
                  --      if txd_rd_pntr is between 0x0 and 0x1F5 then an update of 10 or more words occurred
                    if wrote_first_packet = '0' then
                      set_first_packet <= '1';
                    else
                      set_first_packet <= '0';
                    end if;
                    update_rd_pntrs  <= '0';
                    halt_pntr_update <= '0';
                    disable_txd_trdy <= '0';
                    clr_full_pntr    <= '1';
                    clr_all_hits     <= '1';
                    clr_txd_rdy      <= '0';
                    txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                  else
                  --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                  --    txd_rd_pntr >= txd_rd_pntr_hold
                    update_rd_pntrs  <= '1';
                    halt_pntr_update <= '1';
                    disable_txc_trdy <= '1';
                    disable_txd_trdy <= '1';
                    clr_full_pntr    <= '0';
                    txd_wr_ns        <= CLR_WORDS;
                  end if;
                else
                --  txd_rd_pntr = 0x1F7, 0x1F8, 0x1F9, 0x1FA, 0x1FB, 0x1FC, 0x1FD, 0x1FE, or 0x1FF for 2048 byte memory,
                --  so the minimum txd_rd_pntr_hold_plus9 can be is 0, 1, 2, 3, 4, 5, 6, 7, or 8
                  if (txd_rd_pntr > txd_rd_pntr_hold_plus9) and (txd_rd_pntr < txd_rd_pntr_hold) then
                  --  txd_rd_pntr_hold will be either 0x1F7, 0x1F8, 0x1F9, 0x1FA, 0x1FB, 0x1FC, 0x1FD, 0x1FE, or 0x1FF
                  --  for 2048 byte memory
                  --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                  --      then the update was >= 10 words and the state can be exited
                  --          if  txd_rd_pntr_hold = 0x1F7 then  txd_rd_pntr_hold_plus9 = 0
                  --            txd_rd_pntr has to between 0x1 and 0x1F6 to exit this state
                  --          if  txd_rd_pntr_hold = 0x1F8 then  txd_rd_pntr_hold_plus9 = 1
                  --            txd_rd_pntr has to between 0x2 and 0x1F7 to exit this state
                  --          if  txd_rd_pntr_hold = 0x1F9 then  txd_rd_pntr_hold_plus9 = 2
                  --            txd_rd_pntr has to between 0x3 and 0x1F8 to exit this state
                  --          if  txd_rd_pntr_hold = 0x1FA then  txd_rd_pntr_hold_plus9 = 3
                  --            txd_rd_pntr has to between 0x4 and 0x1F9 to exit this state
                  --          if  txd_rd_pntr_hold = 0x1FB then  txd_rd_pntr_hold_plus9 = 4
                  --            txd_rd_pntr has to between 0x5 and 0x1FA to exit this state
                  --          if  txd_rd_pntr_hold = 0x1FC then  txd_rd_pntr_hold_plus9 = 5
                  --            txd_rd_pntr has to between 0x6 and 0x1FB to exit this state
                  --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus9 = 6
                  --            txd_rd_pntr has to between 0x7 and 0x1FC to exit this state
                  --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus9 = 7
                  --            txd_rd_pntr has to between 0x8 and 0x1FD to exit this state
                  --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus9 = 8
                  --            txd_rd_pntr has to between 0x9 and 0x1FE to exit this state
                    if wrote_first_packet = '0' then
                      set_first_packet <= '1';
                    else
                      set_first_packet <= '0';
                    end if;
                    update_rd_pntrs  <= '0';
                    halt_pntr_update <= '0';
                    disable_txd_trdy <= '0';
                    clr_full_pntr    <= '1';
                    clr_txd_rdy      <= '0';
                    clr_all_hits     <= '1';
                    txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                  else
                  --  txd_rd_pntr did not update by 10 or more words, so update hold poointers and stay in this state
                  --  txd_rd_pntr_hold will be either 0x1F7, 0x1F8, 0x1F9, 0x1FA, 0x1FB, 0x1FC, 0x1FD, 0x1FE, or 0x1FF
                  --  for 2048 byte memory
                  --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                  --      then the update was >= 10 words and the state can be exited BUT
                  --          if  txd_rd_pntr_hold = 0x1F7 then  txd_rd_pntr_hold_plus9 = 0
                  --            txd_rd_pntr was only updated 1-9 words to 0x1F8 - 0x0, so stay here
                  --          if  txd_rd_pntr_hold = 0x1F8 then  txd_rd_pntr_hold_plus9 = 1
                  --            txd_rd_pntr was only updated 1-9 words to 0x1F9 - 0x01 or 0x1, so stay here
                  --          if  txd_rd_pntr_hold = 0x1F9 then  txd_rd_pntr_hold_plus9 = 2
                  --            txd_rd_pntr was only updated 1-9 words to 0x1FA - 0x02 so stay here
                  --          if  txd_rd_pntr_hold = 0x1FA then  txd_rd_pntr_hold_plus9 = 3
                  --            txd_rd_pntr was only updated 1-9 words to 0x1FB - 0x3, so stay here
                  --          if  txd_rd_pntr_hold = 0x1FB then  txd_rd_pntr_hold_plus9 = 4
                  --            txd_rd_pntr was only updated 1-9 words to 0x1FC - 0x4, so stay here
                  --          if  txd_rd_pntr_hold = 0x1FC then  txd_rd_pntr_hold_plus9 = 5
                  --            txd_rd_pntr was only updated 1-9 words to 0x1FD - 0x5, so stay here
                  --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus9 = 6
                  --            txd_rd_pntr was only updated 1-9 words to 0x1FE - 0x6, so stay here
                  --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus9 = 7
                  --            txd_rd_pntr was only updated 1-9 words to 0x1FF - 0x7, so stay here
                  --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus9 = 8
                  --            txd_rd_pntr was only updated 1-9 words to 0x0 - 0x8, so stay here
                    update_rd_pntrs  <= '1';
                    halt_pntr_update <= '1';
                    disable_txc_trdy <= '1';
                    disable_txd_trdy <= '1';
                    clr_full_pntr    <= '0';
                    txd_wr_ns        <= CLR_WORDS;
                  end if;
                end if;
              end if;
            end if;
          else
          --  the update count is > 9 so get out of this state and accept the next packet.
            update_rd_pntrs  <= '0';
            halt_pntr_update <= '0';
            disable_txd_trdy <= '0';
            clr_full_pntr    <= '1';
            clr_all_hits     <= '1';
            clr_txd_rdy      <= '0';
            txd_wr_ns        <= WAIT_COMPARE_CMPLT;
          end if;

        when WAIT_COMPARE_CMPLT =>
          txd_wr_ns        <= IDLE;

        when others =>
          txd_wr_ns <= IDLE;
      end case;
    end process;

    -----------------------------------------------------------------------------
    -- AXI Stream TX Control State Machine Sequencer
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXD_SEQ : process (AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_wr_cs <= IDLE;
        else
          txd_wr_cs <= txd_wr_ns;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    -- Indicator when performing a write to TxD Memory
    --  clear on axi_str_txd_tlast_dly0 = '1'
    -----------------------------------------------------------------------------
    TXD_RDY_INDICATOR : process (AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rdy <= '0';
        else
          if clr_txd_rdy = '1' then
            txd_rdy <= '0';
          elsif set_txd_rdy = '1' then
            txd_rdy <= '1';
          else
            txd_rdy <= txd_rdy;
          end if;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Filter to indicate first packet was written
    --    Needed for full flag
    -----------------------------------------------------------------------------
    FIRST_PACKET_WROTE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          wrote_first_packet     <= '0';
        elsif set_first_packet = '1' then
          wrote_first_packet     <= '1';
        else
          wrote_first_packet     <= wrote_first_packet;
        end if;
      end if;
    end process;

    axi_str_txd_2_mem_addr_int_plus1  <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 1);
    axi_str_txd_2_mem_addr_int_plus3  <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 3);
    axi_str_txd_2_mem_addr_int_plus4  <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 4);
    axi_str_txd_2_mem_addr_int_plus10 <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 10);
    ---------------------------------------------------------------------------
    --  Register to help fmax
    --  With ASYNC BRAM clock cannot read/write same address in memory at same
    --  time unless timing is met, so read until data matches
    ---------------------------------------------------------------------------
    RD_PNTR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rd_pntr_1 <= (others => '0');
          txd_rd_pntr   <= (others => '0');
          compare_addr0_cmplt <= '0';
        else
          if set_txc_addr_0 = '1' and txc_addr_0_dly2 = '1' and
             txc_we_dly2 = '0'  then
          --  txc_addr_0_dly2 is when data is first avaliable from memory

          --  use set_txc_addr_0 to disable compare_addr0_cmplt once pointers update
          --  once state machine advances, set_txc_addr_0 will go low so use it to disable any more
          --  any more data from memory
            txd_rd_pntr_1      <= Axi_Str_TxC_2_Mem_Dout(c_TxD_addrb_width -1 downto 0);

            if Axi_Str_TxC_2_Mem_Dout(c_TxD_addrb_width -1 downto 0) = txd_rd_pntr_1 and
              compare_addr0_cmplt = '0' then
              txd_rd_pntr         <= txd_rd_pntr_1;
              if enable_compare_addr0_cmplt = '1' then
                compare_addr0_cmplt <= '1';
              else
                compare_addr0_cmplt <= '0';
              end if;
            else
              txd_rd_pntr         <= txd_rd_pntr;
              compare_addr0_cmplt <= '0';
            end if;
          else
            txd_rd_pntr_1      <= txd_rd_pntr_1;
            txd_rd_pntr        <= txd_rd_pntr;
            compare_addr0_cmplt<= '0';
          end if;
        end if;
      end if;
    end process;


    ---------------------------------------------------------------------------
    --  Update the read pointer locations until the memory goes FULL
    --    Then use the stored values to compare against real time read pointer
    --    and throttle appropriately
    ---------------------------------------------------------------------------
    RD_PNTRS : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rd_pntr_hold_plus3 <= txc_rd_addr3;
          txd_rd_pntr_hold_plus9 <= txc_rd_addr9;
          txd_rd_pntr_hold       <= txc_rd_addr0;
        else
          if (txd_mem_full = '0' and txc_addr_0_dly2 = '1' and halt_pntr_update = '0') or update_rd_pntrs = '1' then
          --  halt_pntr_update is for the special case when memory is almost full/full and
          --  the Txd FSM needs to wait for a few reads before the next packet starts
          --  The TxD FSM will assert it HIGH to prevent the poiners from being updated
            txd_rd_pntr_hold_plus3 <= std_logic_vector(unsigned(txd_rd_pntr) +3);
            txd_rd_pntr_hold_plus9 <= std_logic_vector(unsigned(txd_rd_pntr) +9);
            txd_rd_pntr_hold       <= txd_rd_pntr;
          else
            txd_rd_pntr_hold_plus3 <= txd_rd_pntr_hold_plus3;
            txd_rd_pntr_hold_plus9 <= txd_rd_pntr_hold_plus9;
            txd_rd_pntr_hold       <= txd_rd_pntr_hold;
          end if;
        end if;
      end if;
    end process;



    ---------------------------------------------------------------------------
    --  Update the read pointer counter to keep ttrack of the total read pointer update is small packets
    --  are sent such that the read pointer is only updated by < 10 words.
    --    This could take up to 4 packets for the read pointer to update to > 10 words
    ---------------------------------------------------------------------------
    RD_PNTR_CNT_UPDATE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
          update_cnt <= (others => '0');
        else
          if update_rd_pntrs = '1' then
            update_cnt <= std_logic_vector(unsigned(update_cnt) + (unsigned(txd_rd_pntr) - unsigned(txd_rd_pntr_hold)));
          else
            update_cnt <= update_cnt;
          end if;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Full flag indicator
    --    Does not begin comparison until 1st packet is written to memory
    -----------------------------------------------------------------------------
    TXD_FULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
            txd_mem_full     <= '0';
            txd_mem_not_full <= '1';
        else
            if (axi_str_txd_2_mem_addr_int_plus3 = txd_rd_pntr and
              (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) then
              txd_mem_full     <= '1';
              txd_mem_not_full <= '0';
            else
              txd_mem_full     <= txd_mem_full;
              txd_mem_not_full <= txd_mem_not_full;
            end if;
        end if;
      end if;
    end process;

    TXD_AFULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
            txd_mem_afull     <= '0';
        else

          if (axi_str_txd_2_mem_addr_int_plus4 = txd_rd_pntr and
              (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) then
            txd_mem_afull     <= '1';
          else
            txd_mem_afull     <= txd_mem_afull;
          end if;
        end if;
      end if;
    end process;


--    TXD_CLR_WORDS_FLAG : process(AXI_STR_TXD_ACLK)
--    begin
--
--      if rising_edge(AXI_STR_TXD_ACLK) then
--        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
--            txd_mem_clr_words     <= '0';
--        else
--
--          if (axi_str_txd_2_mem_addr_int_plus10 = txd_rd_pntr and
--              (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) then
--            txd_mem_clr_words     <= '1';
--          else
--            txd_mem_clr_words     <= txd_mem_clr_words;
--          end if;
--        end if;
--      end if;
--    end process;

    TXD_CLR_WORDS_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
            txd_mem_clr_words     <= '0';
        elsif clr_full_pntr = '1' then
        --  need to take into account if update_cnt <= nine
          if update_cnt <= nine then
          --  once set only clear if conditions are met to allow it to be re-asserted
            if txd_rd_pntr_hold <= txd_max_wr_addr_minus10 then
            --  txd_rd_pntr is between 0x0 and 0x1F5
              if  txd_rd_pntr > txd_rd_pntr_hold_plus9 then              
                -- txd_rd_pntr updated more than 9
                txd_mem_clr_words     <= '0';
              else
                if txd_rd_pntr < txd_rd_pntr_hold then
                --  the read pointer wrapped, so update was greater than 9
                  txd_mem_clr_words     <= '0';  
                else
                  txd_mem_clr_words     <= '1';
                end if;
              end if;
            else
              if txd_rd_pntr_hold_plus9 = txd_max_wr_addr then
              --  txd_rd_pntr = 0x1F6, so any update in which txd_rd_pntr < txd_rd_pntr_hold_plus9
              --  is good
                if txd_rd_pntr <= txd_rd_pntr_hold then
                --  txd_rd_pntr must be 0x0 - 0x1F6
                  txd_mem_clr_words     <= '0';   
                else
                  txd_mem_clr_words     <= '1';
                end if;
              else
                if ((txd_rd_pntr > txd_rd_pntr_hold_plus9) and
                    (txd_rd_pntr < txd_rd_pntr_hold      )) then 
                  txd_mem_clr_words     <= '0';
                else
                  txd_mem_clr_words     <= '1';
                end if;
              end if;
            end if;
          else
            txd_mem_clr_words     <= '0';
          end if;
        else  --set condition

          if (axi_str_txd_2_mem_addr_int_plus10 = txd_rd_pntr and
              (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) then
            txd_mem_clr_words     <= '1';
          else
            txd_mem_clr_words     <= txd_mem_clr_words;
          end if;
        end if;
      end if;
    end process;
    
    
    DELAY_TXD_TREADY_DISABLE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        disable_txd_trdy_dly <= disable_txd_trdy or txd_throttle;
      end if;
    end process;

    DELAY_TREADY_DISABLE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        disable_txc_trdy_dly <= disable_txc_trdy;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  TxD Ready
    --    Only assert when FIFO is not full and TxC is not in process
    -----------------------------------------------------------------------------
    TXD_READY : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_tready_int_dly <= axi_str_txd_tready_int;
        if (AXI_STR_TXD_TLAST = '1' and AXI_STR_TXD_TVALID = '1' and axi_str_txd_tready_int = '1') or
           (clr_txd_trdy = '1' and disable_txd_trdy_dly = '0') or
           disable_txd_trdy = '1' or txd_throttle = '1' then
          axi_str_txd_tready_int <= '0';
        elsif set_txd_rdy = '1' or (txd_rdy = '1' and clr_txd_rdy = '0') then
            if (axi_str_txd_2_mem_addr_int_plus3 = txd_rd_pntr and
               inc_txd_wr_addr = '1') or
               (clr_full_pntr = '0' and txd_mem_full = '1') then
            --  txd_rd_pntr is where the the current read is occuring, so
            --    to account for register pipelines, this needs to stop at
            --    3 counts before the current write address
              axi_str_txd_tready_int <= '0';
            else
              axi_str_txd_tready_int <= '1';
            end if;
        else
          axi_str_txd_tready_int <= '0';
        end if;
      end if;
    end process;

    AXI_STR_TXD_TREADY     <= axi_str_txd_tready_int;


    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_WR_ADDR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_2_mem_addr_int <= (others => '0');
        elsif (inc_txd_wr_addr = '1' or inc_txd_addr_one = '1') then
        --  the address ready for the next transaction
          axi_str_txd_2_mem_addr_int <= std_logic_vector(unsigned(axi_str_txd_2_mem_addr_int) + 1);
        else
          axi_str_txd_2_mem_addr_int <= axi_str_txd_2_mem_addr_int;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Force and update the BRAM with the axi_str_txd_2_mem_addr_int
    --  every ~128 writes (~512 bytes)
    ---------------------------------------------------------------------------
    BRAM_UPDATE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_txd_rdy = '1' then
          update_bram_cnt     <= (others => '0');
        else
          if update_bram_cnt(7) = '1' and inc_txd_wr_addr = '1' then
            update_bram_cnt <= std_logic_vector(unsigned('0' & update_bram_cnt(6 downto 0)) + 1);
          elsif inc_txd_wr_addr = '1' then
            update_bram_cnt <=  std_logic_vector(unsigned(update_bram_cnt) + 1);
          else
            update_bram_cnt <= update_bram_cnt;
          end if;
        end if;
      end if;
    end process;


    axi_str_txd_2_mem_addr               <= axi_str_txd_2_mem_addr_int;


    Axi_Str_TxD_2_Mem_Din(35)           <= axi_str_txd_2_mem_we_int(3);
    Axi_Str_TxD_2_Mem_Din(26)           <= axi_str_txd_2_mem_we_int(2);
    Axi_Str_TxD_2_Mem_Din(17)           <= axi_str_txd_2_mem_we_int(1);
    Axi_Str_TxD_2_Mem_Din(8)            <= axi_str_txd_2_mem_we_int(0);

    Axi_Str_TxD_2_Mem_Din(34 downto 27) <= axi_str_txd_tdata_dly1(31 downto 24);
    Axi_Str_TxD_2_Mem_Din(25 downto 18) <= axi_str_txd_tdata_dly1(23 downto 16);
    Axi_Str_TxD_2_Mem_Din(16 downto  9) <= axi_str_txd_tdata_dly1(15 downto  8);
    Axi_Str_TxD_2_Mem_Din(7  downto  0) <= axi_str_txd_tdata_dly1( 7 downto  0);

    -----------------------------------------------------------------------------
    --  Write Parity bits to the AXI Stream Data Memory
    --    The parity bit always should be the AXI_STR_TXD_TSTRB bits delayed
    -----------------------------------------------------------------------------
    MEM_TXD_PARITY : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_2_mem_we_int <= set_txd_we;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Write Enable bits to the AXI Stream Data Memory
    --    All of the write enables bits should be forced HIGH any time a write to
    --    memory is being performed.  This will allow the parity bits to be
    --    cleared which in turn prevents too much data being read on the Txd
    --    client interface.
    -----------------------------------------------------------------------------
    MEM_TXD_WR_EN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        case set_txd_we is
          when "0000" => Axi_Str_TxD_2_Mem_We <= "0000";
          when others => Axi_Str_TxD_2_Mem_We <= "1111";
        end case;
      end if;
    end process;

--    Axi_Str_TxD_2_Mem_We <= axi_str_txd_2_mem_we_int;

    -----------------------------------------------------------------------------
    --  Enable bit to the AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_EN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if set_txd_en = '1' then
          axi_str_txd_2_mem_en_int <= '1';
        else
          axi_str_txd_2_mem_en_int <= '0';
        end if;
      end if;
    end process;

    Axi_Str_TxD_2_Mem_En <= axi_str_txd_2_mem_en_int;


  -----------------------------------------------------------------------------
  --  VLAN LOGIC
  -----------------------------------------------------------------------------

   ----------------------------------------------------------------------------
   --  Control signal indicating when to check the outter tag for a TPID hit
   ----------------------------------------------------------------------------
   CHECK_TAG0 : process (AXI_STR_TXD_ACLK)
   begin

      if rising_edge(AXI_STR_TXD_ACLK) then
         if setCheckTag0Tpid = '1' then
            checkTag0Tpid <= '1';
         else
            checkTag0Tpid <= '0';
         end if;
         checkTag0Tpid_dly1  <= checkTag0Tpid and not(inhibit_checktag0tpid);
         checkTag0Tpid_dly <= checkTag0Tpid_dly1;
      end if;
   end process;


   ----------------------------------------------------------------------------
   --  Control signal indicating when to check the inner tag for a TPID hit
   ----------------------------------------------------------------------------
   CHECK_TAG1 : process (AXI_STR_TXD_ACLK)
   begin

      if rising_edge(AXI_STR_TXD_ACLK) then
         if setCheckTag1Tpid = '1' then
            checkTag1Tpid <= '1';
         else
            checkTag1Tpid <= '0';
         end if;
         checkTag1Tpid_dly1 <= checkTag1Tpid;
         checkTag1Tpid_dly  <= checkTag1Tpid_dly1;
      end if;
   end process;

   ----------------------------------------------------------------------------
   --  Delay throttle signal
   ----------------------------------------------------------------------------
   DELAY_THROTTLE : process (AXI_STR_TXD_ACLK)
   begin

      if rising_edge(AXI_STR_TXD_ACLK) then
         if txd_throttle = '1' then
            txd_throttle_dly <= '1';
         else
            txd_throttle_dly <= '0';
         end if;
      end if;
   end process;

   ----------------------------------------------------------------------------
   --  Delay throttle signal
   ----------------------------------------------------------------------------
   DELAY_TVALID_IGNORE : process (AXI_STR_TXD_ACLK)
   begin

      if rising_edge(AXI_STR_TXD_ACLK) then
         if ignore_tvalid = '1' then
            ignore_tvalid_dly <= '1';
         else
            ignore_tvalid_dly <= '0';
         end if;
      end if;
   end process;


   ----------------------------------------------------------------------------
   --  Delay throttle signal
   ----------------------------------------------------------------------------
   TXD_TVALID_IGNORE : process (AXI_STR_TXD_ACLK)
   begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_all_hits = '1' then
          ignore_txd_tvalid <= '0';
        else
          if set_ignore_txd_tvalid = '1' then
            ignore_txd_tvalid <= '1';
          else
            ignore_txd_tvalid <= ignore_txd_tvalid;
          end if;
        end if;
      end if;
   end process;


    -----------------------------------------------------------------------------
    --  Enable bit to the Transmit VLAN BRAM
    -----------------------------------------------------------------------------
    TX_VLAN_BRAM_ENABLE : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then -- mw 0510_2011 or clr_vlan_bram_en = '1' then
          tx_vlan_bram_en_int <= '0';
        elsif set_vlan_bram_en = '1' then
          tx_vlan_bram_en_int <= '1';
        else
          tx_vlan_bram_en_int <= '0';--tx_vlan_bram_en_int; --mw 0510_2011
        end if;
        tx_vlan_bram_en_dly1 <= tx_vlan_bram_en_int;
        tx_vlan_bram_en_dly2 <= tx_vlan_bram_en_dly1;
      end if;
    end process;

    tx_vlan_bram_en <= tx_vlan_bram_en_int;
        
    -----------------------------------------------------------------------------
    --  Enable bit to the Transmit VLAN BRAM
    -----------------------------------------------------------------------------
    DECODE_DELAY : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if set_decode_dly = '1' then
          decode_dly1 <= '1';
        else
          decode_dly1 <= '0';
        end if;
        decode_dly2 <= decode_dly1;
        decode_dly3 <= decode_dly2;
        decode_dly4 <= decode_dly3;
        
      end if;
    end process;    
    

    -----------------------------------------------------------------------------
    --  Address to the Transmit VLAN BRAM
    -----------------------------------------------------------------------------
    TX_VLAN_BRAM_ADDRESS : process(tx_vlan_bram_en_int,axi_str_txd_tdata_dly0)
    begin
      if tx_vlan_bram_en_int = '1' then
        tx_vlan_bram_addr_int <= axi_str_txd_tdata_dly0(19 downto 16) & axi_str_txd_tdata_dly0(31 downto 24);
      else
        tx_vlan_bram_addr_int <= (others => '0');
      end if;
    end process;

    tx_vlan_bram_addr <= tx_vlan_bram_addr_int;

    REG_BRAM_DIN : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if tx_vlan_bram_en_dly1 = '1' then
          tx_vlan_bram_din_dly <= tx_vlan_bram_din;
        else
          tx_vlan_bram_din_dly <= (others => '0');
        end if;
      end if;
    end process;

end rtl;


-------------------------------------------------------------------------------
-- tx_csum_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_csum_if.vhd
-- Version:         v1.00a
-- Description:     top level of embedded ip Ethernet MAC interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--                    tx_axistream_if.vhd
--          ->          tx_csum_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd

--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

library work;
use work.tx_if_pack.all;



-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity tx_csum_if is
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0)   --  Tx AXI-Stream Control to Memory Full Flag

  );

end tx_csum_if;
------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of tx_csum_if is
begin

-------------------------------------------------------------------------------
--  Start Partial CSUM
-------------------------------------------------------------------------------
GEN_CSUM_PARTIAL : if (C_TXCSUM  = 1 and (C_TXVLAN_TRAN = 0 and C_TXVLAN_TAG = 0 and C_TXVLAN_STRP = 0)) generate
begin

  TX_CSUM_PARTIAL_INTERFACE : tx_csum_partial_if
  --  Interface for Transmit AxiStream Data and Control; and Tx Memory
  generic map (
    C_FAMILY               => C_FAMILY,
    C_HALFDUP              => C_HALFDUP,
    C_TXCSUM               => C_TXCSUM,
    C_TXMEM                => C_TXMEM,
    C_TXVLAN_TRAN          => C_TXVLAN_TRAN,
    C_TXVLAN_TAG           => C_TXVLAN_TAG,
    C_TXVLAN_STRP          => C_TXVLAN_STRP,
    C_S_AXI_ADDR_WIDTH     => C_S_AXI_ADDR_WIDTH,
    C_S_AXI_DATA_WIDTH     => C_S_AXI_DATA_WIDTH,

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    => c_TxD_write_width_b,
    c_TxD_read_width_b     => c_TxD_read_width_b,
    c_TxD_write_depth_b    => c_TxD_write_depth_b,
    c_TxD_read_depth_b     => c_TxD_read_depth_b,
    c_TxD_addrb_width      => c_TxD_addrb_width,
    c_TxD_web_width        => c_TxD_web_width,

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    => c_TxC_write_width_b,
    c_TxC_read_width_b     => c_TxC_read_width_b,
    c_TxC_write_depth_b    => c_TxC_write_depth_b,
    c_TxC_read_depth_b     => c_TxC_read_depth_b,
    c_TxC_addrb_width      => c_TxC_addrb_width,
    c_TxC_web_width        => c_TxC_web_width

  )
  port map  (

    tx_init_in_prog        => tx_init_in_prog,

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       => AXI_STR_TXD_ACLK,
    reset2axi_str_txd      => reset2axi_str_txd,
    AXI_STR_TXD_TVALID     => AXI_STR_TXD_TVALID,
    AXI_STR_TXD_TREADY     => AXI_STR_TXD_TREADY,
    AXI_STR_TXD_TLAST      => AXI_STR_TXD_TLAST,
    AXI_STR_TXD_TSTRB      => AXI_STR_TXD_TSTRB,
    AXI_STR_TXD_TDATA      => AXI_STR_TXD_TDATA,
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       => AXI_STR_TXC_ACLK,
    reset2axi_str_txc      => reset2axi_str_txc,
    AXI_STR_TXC_TVALID     => AXI_STR_TXC_TVALID,
    AXI_STR_TXC_TREADY     => AXI_STR_TXC_TREADY,
    AXI_STR_TXC_TLAST      => AXI_STR_TXC_TLAST,
    AXI_STR_TXC_TSTRB      => AXI_STR_TXC_TSTRB,
    AXI_STR_TXC_TDATA      => AXI_STR_TXC_TDATA,

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  => Axi_Str_TxD_2_Mem_Din,       --: out std_logic_vector(c_TxD_write_width_b-1 downto 0);
    Axi_Str_TxD_2_Mem_Addr => Axi_Str_TxD_2_Mem_Addr,      --: out std_logic_vector(c_TxD_addrb_width-1   downto 0);
    Axi_Str_TxD_2_Mem_En   => Axi_Str_TxD_2_Mem_En,        --: out std_logic := '1';
    Axi_Str_TxD_2_Mem_We   => Axi_Str_TxD_2_Mem_We,        --: out std_logic_vector(c_TxD_web_width-1     downto 0);
    Axi_Str_TxD_2_Mem_Dout => Axi_Str_TxD_2_Mem_Dout,      --: in  std_logic_vector(c_TxD_read_width_b-1  downto 0);

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  => Axi_Str_TxC_2_Mem_Din,       --: out std_logic_vector(c_TxD_write_width_b-1 downto 0);
    Axi_Str_TxC_2_Mem_Addr => Axi_Str_TxC_2_Mem_Addr,      --: out std_logic_vector(c_TxD_addrb_width-1   downto 0);
    Axi_Str_TxC_2_Mem_En   => Axi_Str_TxC_2_Mem_En,        --: out std_logic := '1';
    Axi_Str_TxC_2_Mem_We   => Axi_Str_TxC_2_Mem_We,        --: out std_logic_vector(c_TxD_web_width-1     downto 0);
    Axi_Str_TxC_2_Mem_Dout => Axi_Str_TxC_2_Mem_Dout       --: in  std_logic_vector(c_TxD_read_width_b-1  downto 0);

  );
end generate GEN_CSUM_PARTIAL;
-------------------------------------------------------------------------------
--  End Partial CSUM
-------------------------------------------------------------------------------


-------------------------------------------------------------------------------
--  Start FULL CSUM
-------------------------------------------------------------------------------
GEN_CSUM_FULL : if (C_TXCSUM  = 2 and (C_TXVLAN_TRAN = 0 and C_TXVLAN_TAG = 0 and C_TXVLAN_STRP = 0)) generate
begin

  TX_CSUM_FULL_INTERFACE : tx_csum_full_if
  --  Interface for Transmit AxiStream Data and Control; and Tx Memory
  generic map (
    C_FAMILY               => C_FAMILY,
    C_HALFDUP              => C_HALFDUP,
    C_TXCSUM               => C_TXCSUM,
    C_TXMEM                => C_TXMEM,
    C_TXVLAN_TRAN          => C_TXVLAN_TRAN,
    C_TXVLAN_TAG           => C_TXVLAN_TAG,
    C_TXVLAN_STRP          => C_TXVLAN_STRP,
    C_S_AXI_ADDR_WIDTH     => C_S_AXI_ADDR_WIDTH,
    C_S_AXI_DATA_WIDTH     => C_S_AXI_DATA_WIDTH,

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    => c_TxD_write_width_b,
    c_TxD_read_width_b     => c_TxD_read_width_b,
    c_TxD_write_depth_b    => c_TxD_write_depth_b,
    c_TxD_read_depth_b     => c_TxD_read_depth_b,
    c_TxD_addrb_width      => c_TxD_addrb_width,
    c_TxD_web_width        => c_TxD_web_width,

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    => c_TxC_write_width_b,
    c_TxC_read_width_b     => c_TxC_read_width_b,
    c_TxC_write_depth_b    => c_TxC_write_depth_b,
    c_TxC_read_depth_b     => c_TxC_read_depth_b,
    c_TxC_addrb_width      => c_TxC_addrb_width,
    c_TxC_web_width        => c_TxC_web_width

  )
  port map  (

    tx_init_in_prog        => tx_init_in_prog,

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       => AXI_STR_TXD_ACLK,
    reset2axi_str_txd      => reset2axi_str_txd,
    AXI_STR_TXD_TVALID     => AXI_STR_TXD_TVALID,
    AXI_STR_TXD_TREADY     => AXI_STR_TXD_TREADY,
    AXI_STR_TXD_TLAST      => AXI_STR_TXD_TLAST,
    AXI_STR_TXD_TSTRB      => AXI_STR_TXD_TSTRB,
    AXI_STR_TXD_TDATA      => AXI_STR_TXD_TDATA,
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       => AXI_STR_TXC_ACLK,
    reset2axi_str_txc      => reset2axi_str_txc,
    AXI_STR_TXC_TVALID     => AXI_STR_TXC_TVALID,
    AXI_STR_TXC_TREADY     => AXI_STR_TXC_TREADY,
    AXI_STR_TXC_TLAST      => AXI_STR_TXC_TLAST,
    AXI_STR_TXC_TSTRB      => AXI_STR_TXC_TSTRB,
    AXI_STR_TXC_TDATA      => AXI_STR_TXC_TDATA,

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  => Axi_Str_TxD_2_Mem_Din,       --: out std_logic_vector(c_TxD_write_width_b-1 downto 0);
    Axi_Str_TxD_2_Mem_Addr => Axi_Str_TxD_2_Mem_Addr,      --: out std_logic_vector(c_TxD_addrb_width-1   downto 0);
    Axi_Str_TxD_2_Mem_En   => Axi_Str_TxD_2_Mem_En,        --: out std_logic := '1';
    Axi_Str_TxD_2_Mem_We   => Axi_Str_TxD_2_Mem_We,        --: out std_logic_vector(c_TxD_web_width-1     downto 0);
    Axi_Str_TxD_2_Mem_Dout => Axi_Str_TxD_2_Mem_Dout,      --: in  std_logic_vector(c_TxD_read_width_b-1  downto 0);

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  => Axi_Str_TxC_2_Mem_Din,       --: out std_logic_vector(c_TxD_write_width_b-1 downto 0);
    Axi_Str_TxC_2_Mem_Addr => Axi_Str_TxC_2_Mem_Addr,      --: out std_logic_vector(c_TxD_addrb_width-1   downto 0);
    Axi_Str_TxC_2_Mem_En   => Axi_Str_TxC_2_Mem_En,        --: out std_logic := '1';
    Axi_Str_TxC_2_Mem_We   => Axi_Str_TxC_2_Mem_We,        --: out std_logic_vector(c_TxD_web_width-1     downto 0);
    Axi_Str_TxC_2_Mem_Dout => Axi_Str_TxC_2_Mem_Dout       --: in  std_logic_vector(c_TxD_read_width_b-1  downto 0);

  );
end generate GEN_CSUM_FULL;
-------------------------------------------------------------------------------
--  End FULL CSUM
-------------------------------------------------------------------------------


end rtl;


-------------------------------------------------------------------------------
-- tx_basic_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_basic_if.vhd
-- Version:         v1.00a
-- Description:     embedded ip AXI Stream transmit interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--                    tx_axistream_if.vhd
--          ->          tx_basic_if.vhd
--                      tx_csum_if.vhd
--                        tx_csum_partial_if.vhd
--                          tx_csum_partial_calc_if.vhd
--                        tx_full_csum_if.vhd
--                      tx_vlan_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tx_if_pack.all;

-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity tx_basic_if is
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    tx_init_in_prog        : out std_logic;                                         --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                         --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                         --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                         --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                         --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                         --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                         --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);   --  AXI-Stream Transmit Control Data

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);  --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);  --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);  --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);  --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                         --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);  --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0)   --  Tx AXI-Stream Control to Memory Full Flag

  );

end tx_basic_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of tx_basic_if is

-------------------------------------------------------------------------------
--  Start Basic Design - No CSUM,  No Extended VLAN
-------------------------------------------------------------------------------

  constant zeroes_txc    : std_logic_vector(c_TxC_write_width_b -1 downto c_TxC_addrb_width) := (others => '0');
  constant zeroes_txd    : std_logic_vector(c_TxC_write_width_b -1 downto c_TxD_addrb_width) := (others => '0');
  constant zeroes_txd_2  : std_logic_vector(c_TxC_write_width_b -1 downto c_TxD_addrb_width + 2 ) := (others => '0');

  type TXC_WR_FSM_TYPE is (
                       TXC_ADDR2_WR,
                       TXC_ADDR0_WR,
                       WAIT_WR_CMPLT,
                       TXC_WD0,
--                       WAIT_TXD_FULL,
                       TXC_WD1,
                       WAIT_ADDR2_COMPARE_CMPLT,--added for BRAM async clocks
                       TXC_WD2,
                       TXC_WD3,
                       TXC_WD4,
                       WAIT_ADDR0_COMPARE_CMPLT,--added for BRAM async clocks
                       TXC_WD5,
                       WAIT_TXD_CMPLT,
                       WAIT_TXD_MEM,
                       WR_TXC_PNTR,
                       WR_TXD_END_PNTR
                      );
  signal txc_wr_cs, txc_wr_ns             : TXC_WR_FSM_TYPE;

  type TXD_WR_FSM_TYPE is (
                       IDLE,
                       TXD_PRM,
                       TXD_WRT,
                       MEM_FULL,
                       CLR_FULL,
                       WAIT_WR1,
                       WAIT_WR2,
                       WAIT_COMPARE_CMPLT
                      );
  signal txd_wr_cs, txd_wr_ns             : TXD_WR_FSM_TYPE;

  signal txc_min_wr_addr                  : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_rsvd_wr_addr                 : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_max_wr_addr                  : std_logic_vector(c_TxC_addrb_width -1 downto 0);

  signal txc_wr_addr0                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr1                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr2                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr3                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr5                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);
  signal txc_wr_addr6                     : std_logic_vector(c_TxC_addrb_width -1 downto 0);

  signal axi_str_txc_tready_int           : std_logic;
  signal axi_str_txc_tready_int_dly       : std_logic;
  signal axi_str_txc_tvalid_dly0          : std_logic;
  signal axi_str_txc_tlast_dly0           : std_logic;
--  signal axi_str_txc_tstrb_dly0           : std_logic_vector(3 downto 0);
  signal axi_str_txc_tdata_dly0           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal clr_txc_trdy                     : std_logic;

  signal axi_str_txd_tready_int           : std_logic;
  signal axi_str_txd_tready_int_dly       : std_logic;
  signal axi_str_txd_tvalid_dly0          : std_logic;
  signal axi_str_txd_tlast_dly0           : std_logic;
  signal axi_str_txd_tstrb_dly0           : std_logic_vector(3 downto 0);
  signal axi_str_txd_tdata_dly0           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal axi_str_txd_tdata_dly1           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
  signal clr_txd_trdy                     : std_logic;

  signal set_txc_addr_0                   : std_logic;
  signal txc_addr_0_dly1                  : std_logic;
  signal txc_addr_0_dly2                  : std_logic;
  signal set_txc_addr_1                   : std_logic;
  signal txc_addr_1                       : std_logic;
  signal set_txc_addr_2                   : std_logic;
  signal txc_addr_2                       : std_logic;
  signal set_txc_addr_4_n                 : std_logic;
  signal set_txc_addr_3                   : std_logic;
  signal clr_txc_addr_3                   : std_logic;
  signal txc_addr_3_dly                   : std_logic;
  signal txc_addr_3_dly2                  : std_logic;
  signal txc_addr_3_dly3                  : std_logic;
  signal inc_txd_addr_one                 : std_logic;
  signal set_txc_trdy                     : std_logic;
  signal set_txc_trdy2                    : std_logic;
  signal clr_txc_trdy2                    : std_logic;
  signal set_txcwr_rd_addr                : std_logic;
  signal set_txcwr_wr_end                 : std_logic;
  signal set_txc_en                       : std_logic;
  signal set_txc_we                       : std_logic;
  signal txc_we                           : std_logic;
  signal txc_we_dly1                      : std_logic;
  signal txc_we_dly2                      : std_logic;
  signal addr_2_en                        : std_logic;
  signal addr_2_en_dly1                   : std_logic;
  signal addr_2_en_dly2                   : std_logic;

  signal txc_mem_full                     : std_logic;
  signal txc_mem_not_full                 : std_logic;
  signal txc_mem_afull                    : std_logic;
  signal txc_mem_wr_addr                  : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_0                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_1                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_last             : std_logic_vector(c_TxC_addrb_width   -1 downto 0);

  signal Axi_Str_TxC_2_Mem_Addr_int       : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal Axi_Str_TxC_2_Mem_We_int         : std_logic_vector(0 downto 0);
  signal txc_mem_wr_addr_plus1            : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_mem_wr_addr_plus2            : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_rd_addr2_pntr                : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal txc_rd_addr2_pntr_1              : std_logic_vector(c_TxC_addrb_width   -1 downto 0);


  -- Set to the full width of the write data bus
  signal Axi_Str_TxC_2_Mem_Din_int        : std_logic_vector(c_TxC_write_width_b -1 downto 0);

  signal set_axi_flag                     : std_logic;
  signal set_csum_cntrl                   : std_logic;
  signal set_csum_begin_insert            : std_logic;
  signal set_csum_rsvd_init               : std_logic;
  signal axi_flag                         : std_logic_vector( 3 downto 0);
  signal csum_cntrl                       : std_logic_vector( 1 downto 0);

  signal set_first_packet                 : std_logic;
  signal wrote_first_packet               : std_logic;
  signal inc_txd_wr_addr                  : std_logic;
  signal set_txd_we                       : std_logic_vector( 3 downto 0);
  signal set_txd_en                       : std_logic;
  signal set_txd_rdy                      : std_logic;
  signal clr_txd_rdy                      : std_logic;
  signal clr_full_pntr                    : std_logic;
  signal halt_pntr_update                 : std_logic;
  signal disable_txd_trdy                 : std_logic;
  signal disable_txd_trdy_dly             : std_logic;
  signal disable_txc_trdy                 : std_logic;
  signal disable_txc_trdy_dly             : std_logic;

  signal txd_rdy                          : std_logic;
  signal axi_str_txd_2_mem_addr_int       : unsigned(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus1 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus2 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus3 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal axi_str_txd_2_mem_addr_int_plus4 : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txd_mem_full                     : std_logic;
  signal txd_mem_not_full                 : std_logic;
  signal txd_mem_afull                    : std_logic;
  signal axi_str_txd_2_mem_we_int         : std_logic_vector( 3 downto 0);
  signal axi_str_txd_2_mem_en_int         : std_logic;

  signal txd_rd_pntr                      : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_1                    : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_reg                  : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_min_wr_addr                  : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_max_wr_addr                  : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_max_wr_addr_minus4           : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_hold_plus3           : std_logic_vector(c_TxD_addrb_width -1 downto 0);
  signal txd_rd_pntr_hold                 : std_logic_vector(c_TxD_addrb_width -1 downto 0);

  signal tx_init_in_prog_int              : std_logic;
  signal init_bram                        : std_logic;

  signal txc_rd_addr0                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txc_rd_addr2                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal txc_rd_addr3                     : std_logic_vector(c_TxD_addrb_width   -1 downto 0);


  signal compare_addr0                    : std_logic;
  signal compare_addr0_cmplt              : std_logic;

  signal compare_addr2                    : std_logic;
  signal compare_addr2_cmplt              : std_logic;
  signal compare_addr2_cmplt_dly          : std_logic;

  signal update_bram_cnt                  : std_logic_vector(7 downto 0);

  signal enable_compare_addr0_cmplt       : std_logic;
  signal end_addr_byte_offset             : std_logic_vector(1 downto 0);
  signal check_full                       : std_logic;
  signal update_rd_pntrs                  : std_logic;

  begin

    -----------------------------------------------------------------------------
    --  The TxC BRAM is set up to to always store the current TxD Read and Write
    --    pointers in the first two locations (0x0 and 0x1) of the Memory
    --    respectivively.  The current TxC Read and write pointer are always
    --    stored in the the next two locations (0x2 and 0x3) of the Memory
    --    respectively.  The End addresses for each packet are then stored
    --    in the remaing Memory locations starting at address 0x4.  After
    --    the end pointer to the maximum address has been written, if the
    --    memory is not full, the address pointer will loop back to address
    --    0x4 and write the end pointer for the next packet.
    --
    --                                   BRAM
    --                             Write       Read
    --                           _____________________
    --                          |__________|_________| <-- TxD Rd Pointer
    --      TxD Wr Pointer -->  |__________|_________|
    --                          |__________|_________| <-- TxC Rd Pointer
    --      TxC Wr Pointer -->  |__________|_________|
    --      Packet 0 End   -->  |__________|_________|  --> Packet 0 End
    --      Packet 1 End   -->  |__________|_________|  --> Packet 1 End
    --      Packet 2 End   -->  |__________|_________|  --> Packet 2 End
    --         .                |__________|_________|         .
    --         .                |__________|_________|         .
    --         .                |__________|_________|         .
    --      Packet n End   -->  |__________|_________|  --> Packet n End
    --
    -----------------------------------------------------------------------------

    -----------------------------------------------------------------------------
    --  Create the full and empty comparison values for the S6 and V6 since
    --  1 S6 BRAM = 1/2 V6 BRAM
    -----------------------------------------------------------------------------
    GEN_TXC_MIN_MAX_WR_FLAG : for i in (c_TxC_addrb_width-1) downto 0 generate
      txc_min_wr_addr(i)  <= '1' when (i = 2)          else '0'; -- do not loop back to 0x0; loop to 0x4
      txc_max_wr_addr(i)  <= '0' when (i = 0 or i = 1) else '1';
      txc_wr_addr0(i)     <= '0';
      txc_wr_addr1(i)     <= '1' when (i = 0)          else '0';
      txc_wr_addr2(i)     <= '1' when (i = 1)          else '0';
      txc_wr_addr3(i)     <= '1' when (i = 0 or i = 1) else '0';
      txc_wr_addr5(i)     <= '1' when (i = 0 or i = 2) else '0';
      txc_wr_addr6(i)     <= '1' when (i = 1 or i = 2) else '0';
    end generate GEN_TXC_MIN_MAX_WR_FLAG;

    GEN_TXD_MIN_MAX_WR_FLAG : for i in (c_TxD_addrb_width-1) downto 0 generate
      txd_min_wr_addr(i)        <= '1' when (i = 0) else '0';
      txd_max_wr_addr_minus4(i) <= '0' when (i = 2) else '1';
      txd_max_wr_addr(i)        <= '1';
    end generate GEN_TXD_MIN_MAX_WR_FLAG;


    GEN_TXC_MIN_MAX_RD_FLAG : for i in (c_TxD_addrb_width-1) downto 0 generate
      txc_rd_addr0(i)     <= '0';
      txc_rd_addr2(i)     <= '1' when (i = 1)          else '0';
      txc_rd_addr3(i)     <= '1' when (i = 0 or i = 1) else '0';
    end generate GEN_TXC_MIN_MAX_RD_FLAG;




    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Control Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXC_CONTROL : process(AXI_STR_TXC_ACLK)
    begin
      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          axi_str_txc_tvalid_dly0 <= '0';
          axi_str_txc_tlast_dly0  <= '0';
          clr_txc_trdy           <= '0';
        else
          axi_str_txc_tvalid_dly0 <= axi_str_txc_tvalid;
          axi_str_txc_tlast_dly0  <= axi_str_txc_tlast;
          if axi_str_txc_tvalid = '1' and axi_str_txc_tlast = '1' and axi_str_txc_tready_int = '1' then
            clr_txc_trdy <= '1';
          else
            clr_txc_trdy <= '0';
          end if;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Control Data Bus
    -----------------------------------------------------------------------------
    REG_TXC_IN : process(AXI_STR_TXC_ACLK)
    begin
      if rising_edge(AXI_STR_TXC_ACLK) then
--          axi_str_txc_tstrb_dly0  <= axi_str_txc_tstrb;
          axi_str_txc_tdata_dly0  <= axi_str_txc_tdata;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  AXI Stream TX Control State Machine - combinational/combinatorial
    --    Used to register the incoming control and checksum information
    --    This state machine will throttle the Transmit AXI Stream Data state
    --      machine until after the control information has been received.
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXC_CMB : process (txc_wr_cs,axi_str_txc_tvalid_dly0,
      axi_str_txc_tlast_dly0,axi_str_txd_tlast_dly0,
      axi_str_txd_tvalid_dly0,txc_addr_3_dly,
      wrote_first_packet,axi_str_txc_tready_int_dly,axi_str_txd_tready_int_dly,
      disable_txd_trdy_dly,disable_txc_trdy_dly,
      compare_addr2_cmplt,compare_addr2_cmplt_dly,compare_addr0_cmplt,
      update_bram_cnt,txc_mem_full)

    begin


      set_axi_flag           <= '0';
      set_csum_cntrl         <= '0';
      set_csum_begin_insert  <= '0';
      set_csum_rsvd_init     <= '0';
      set_txc_addr_0         <= '0';
      set_txc_addr_1         <= '0';
      set_txc_addr_2         <= '0';
      set_txc_addr_3         <= '0';
      set_txc_addr_4_n       <= '0';
      clr_txc_addr_3         <= '0';
      set_txcwr_rd_addr      <= '0';  --  sets the write side, read address to 0x0
      set_txcwr_wr_end       <= '0';  --  writes the end address to the memory in the next available location
      set_txc_en             <= '0';  --  the enable bit to the write side of the memory
      set_txc_we             <= '0';  --  the write enable bit to the write side of the memory
      inc_txd_addr_one       <= '0';
      set_txc_trdy           <= '0';
      init_bram              <= '0';
      compare_addr2          <= '0';
      compare_addr0          <= '0';
      set_txc_trdy2          <= '0';
      clr_txc_trdy2          <= '0';
      enable_compare_addr0_cmplt <= '0';

      case txc_wr_cs is
        when TXC_ADDR2_WR =>
          set_txc_addr_2         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          txc_wr_ns              <= TXC_ADDR0_WR;
        when TXC_ADDR0_WR =>
          set_txc_addr_0         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          txc_wr_ns              <= WAIT_WR_CMPLT;
        when WAIT_WR_CMPLT =>
          set_txc_addr_0         <= '1';
          set_txc_en             <= '1';
          set_txc_we             <= '1';
          init_bram              <= '1';
          set_txc_trdy2          <= '1';
          txc_wr_ns              <= TXC_WD0;
        when TXC_WD0 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' and
             (wrote_first_packet = '0' or txc_addr_3_dly = '1') then
            set_txc_addr_2         <= '1';  --Set the address to get the TxC Rd Address Pointer
            set_txc_en             <= '1';
            set_axi_flag           <= '1';
            clr_txc_addr_3         <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD1;
          else
            set_txc_addr_2         <= '0';  --Set the address to get the TxC Rd Address Pointer
            set_txc_en             <= '0';
            set_axi_flag           <= '0';
            clr_txc_addr_3         <= '0';
            compare_addr2          <= '0';
            txc_wr_ns              <= TXC_WD0;
          end if;

        when TXC_WD1 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_txc_trdy2          <= '0';
            set_csum_cntrl         <= '1';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD2;--WAIT_ADDR2_COMPARE_CMPLT;
          elsif axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '0' then
          -- need to force txc trdy HIGH since TVALID throttled
            set_txc_trdy2          <= '1';
            set_csum_cntrl         <= '0';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= WAIT_ADDR2_COMPARE_CMPLT;
          else
            set_txc_trdy2          <= '0';
            set_csum_cntrl         <= '0';
            set_txc_addr_2         <= '1';
            set_txc_en             <= '1';
            compare_addr2          <= '1';
            txc_wr_ns              <= TXC_WD1;
          end if;

        when WAIT_ADDR2_COMPARE_CMPLT =>
        -- now clear txc trdy to only allow a one clock pulse HIGH
          clr_txc_trdy2          <= '1';
          set_txc_addr_2         <= '1';
          set_txc_en             <= '1';
          compare_addr2          <= '1';
          txc_wr_ns              <= TXC_WD1;

        when TXC_WD2 =>
        -- Txc Tready has already been disabled
        --  wait for compare_addr2_cmplt, then
        --  set_txc_trdy2 will force axi_str_txc_tready_int_dly HIGH
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_csum_begin_insert      <= '1';
            set_txc_addr_2         <= '0';
            set_txc_en             <= '0';
            compare_addr2          <= '0';
            set_txc_trdy2          <= '0';
            txc_wr_ns                  <= TXC_WD3;
          else
            if axi_str_txc_tvalid_dly0 = '0'  or
               (txc_mem_full = '1' and axi_str_txc_tvalid_dly0 = '1') then
            --  If full wait for FULL and TVALID
            --  This will allow next elsif to be hit properly
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '1';
              set_txc_en             <= '1';
              compare_addr2          <= '1';
              set_txc_trdy2          <= '0';
              txc_wr_ns              <= TXC_WD2;


            elsif axi_str_txc_tvalid_dly0 = '1' and
              (compare_addr2_cmplt = '1' or compare_addr2_cmplt_dly = '1') then
              --  when full is '0', only need compare_addr2_cmplt to set set_txc_trdy2
              --    which will then allow this state to be exited to TXD_WD3
              --  when full is '1', then will need compare_addr2_cmplt_dly to to set set_txc_trdy2
              --    which will then allow this state to be exited to TXD_WD3
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '0';
              set_txc_en             <= '0';
              compare_addr2          <= '0';
              set_txc_trdy2          <= '1';
              txc_wr_ns                  <= TXC_WD2;
            else
              set_csum_begin_insert  <= '0';
              set_txc_addr_2         <= '1';
              set_txc_en             <= '1';
              compare_addr2          <= '1';
              set_txc_trdy2          <= '0';
              txc_wr_ns                  <= TXC_WD2;
            end if;
          end if;
        when TXC_WD3 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
          --  This is the earliest state to check for TxC FULL from TXC_WD0 state addr_2
          --  Register data, then assert full = 2 clks from rd
          --    Not FULL so write TxC Write Pointer to addr 0x3
            set_csum_rsvd_init         <= '1';
            txc_wr_ns                  <= TXC_WD4;
          else
            set_csum_rsvd_init         <= '0';
            txc_wr_ns                  <= TXC_WD3;
          end if;
        when TXC_WD4 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' then
            set_txc_addr_0             <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            txc_wr_ns                  <= TXC_WD5;
          else
            set_txc_addr_0             <= '0';  --Set the address to get the TxD Rd Address Pointer
            set_txc_en                 <= '0';
            compare_addr0              <= '0';
            txc_wr_ns                  <= TXC_WD4;
          end if;
        when TXC_WD5 =>
          if axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1' and axi_str_txc_tlast_dly0 = '1' then
            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '1';
            txc_wr_ns                  <= WAIT_ADDR0_COMPARE_CMPLT;
          else
            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '0';
            txc_wr_ns                  <= TXC_WD5;
          end if;
        when WAIT_ADDR0_COMPARE_CMPLT =>
          if compare_addr0_cmplt = '1' then
            set_txc_addr_1             <= '1'; -- this is one clock early, so do not set the we enable yet
            set_txc_en                 <= '1';
            set_txc_we                 <= '1';

            set_txc_addr_0             <= '0';
            set_txc_en                 <= '0';
            compare_addr0              <= '0';
            enable_compare_addr0_cmplt <= '0';
            txc_wr_ns                  <= WAIT_TXD_CMPLT;
          else
            set_txc_addr_1             <= '0';
            set_txc_en                 <= '0';
            set_txc_we                 <= '0';

            set_txc_addr_0             <= '1';
            set_txc_en                 <= '1';
            compare_addr0              <= '1';
            enable_compare_addr0_cmplt <= '1';
            txc_wr_ns                  <= WAIT_ADDR0_COMPARE_CMPLT;
          end if;



        when WAIT_TXD_CMPLT =>
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1'  and
             axi_str_txd_tlast_dly0 = '1' then
            set_txc_addr_0        <= '0';
            set_txc_addr_1        <= '1';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WR_TXD_END_PNTR;
          elsif disable_txd_trdy_dly = '1' then
          -- Txd mem is full so get the current read pointer
          --  This can occure after tlast so check it in the following states
            set_txc_addr_0        <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_addr_1        <= '0';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_MEM;
          elsif update_bram_cnt(7) = '1'  then
          --Writing the current TxC write pointer so the read side can monitor it
            set_txc_addr_1        <= '1';
            set_txc_addr_2        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          else
            set_txc_addr_1        <= '0'; --Writing the current TxC write pointer so the read side can monitor it
            set_txc_addr_2        <= '0';
            set_txc_en            <= '0';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          end if;
        when WAIT_TXD_MEM =>
          if disable_txd_trdy_dly = '1' then
            -- Txd mem is full so get the current read pointer
            set_txc_addr_0        <= '1';  --Set the address to get the TxD Rd Address Pointer
            set_txc_addr_1        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            txc_wr_ns             <= WAIT_TXD_MEM;
          else
            set_txc_addr_0        <= '0';
            set_txc_addr_1        <= '1'; -- this is one clock early, so do not set the we enable yet
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WAIT_TXD_CMPLT;
          end if;
        when WR_TXD_END_PNTR =>
            inc_txd_addr_one      <= '1';
            set_txc_addr_4_n      <= '1'; -- Write the TxC End Value to address 0x4 - 0xn
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            txc_wr_ns             <= WR_TXC_PNTR;

        when WR_TXC_PNTR =>
          if disable_txc_trdy_dly = '1' then
            set_txc_addr_0        <= '1';
            set_txc_addr_3        <= '0';
            set_txc_en            <= '1';
            set_txc_we            <= '0';
            set_txc_trdy          <= '0';
            txc_wr_ns             <= WR_TXC_PNTR;
          else
            set_txc_addr_0        <= '0'; -- Write the TxC end pointer value to start the tx clint FSM
            set_txc_addr_3        <= '1';
            set_txc_en            <= '1';
            set_txc_we            <= '1';
            set_txc_trdy          <= '1';
            txc_wr_ns             <= TXC_WD0;
          end if;

--        when WR_TXC_PNTR =>
--            set_txc_addr_3        <= '1'; -- Write the TxC end pointer value to start the tx clint FSM
--            set_txc_addr_0        <= '0';
--            set_txc_en            <= '1';
--            set_txc_we            <= '1';
--            txc_wr_ns             <= TXC_WD0;

        when others =>
          txc_wr_ns                <= TXC_ADDR2_WR;
      end case;
    end process;

    -----------------------------------------------------------------------------
    -- AXI Stream TX Control State Machine Sequencer
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXC_SEQ : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_wr_cs <= TXC_ADDR2_WR;
        else
          txc_wr_cs <= txc_wr_ns;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    -- Delay the last write to TxC memory of the first packet after reset
    -----------------------------------------------------------------------------
    TX_INIT_INDICATOR_DLYS : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_addr_3_dly2 <= '0';
          txc_addr_3_dly3 <= '0';
        else
          txc_addr_3_dly2 <= txc_addr_3_dly;
          txc_addr_3_dly3 <= txc_addr_3_dly2;
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    -- Use above delay to hold off Tx Client FSM from starting until all
    --    TxD and TxC pointer information has been written to memory
    --
    --    This signal goes through a clock crossing circuit before it is
    --      registered in the Tx Client clock domain and used to start the
    --      Tx Client Read FSM
    -----------------------------------------------------------------------------
    TX_INIT_INDICATOR : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          tx_init_in_prog_int <= '1';
        else
          if txc_addr_3_dly3 = '1' then
            tx_init_in_prog_int <= '0';
          else
            tx_init_in_prog_int <= tx_init_in_prog_int;
          end if;
        end if;
      end if;
    end process;

    tx_init_in_prog <= tx_init_in_prog_int;

    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_1_TXD_WR_PNTR : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_1 = '1' then
          txc_addr_1 <= '1';
        else
          txc_addr_1 <= '0';
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_3_DELAY : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' or clr_txc_addr_3 = '1' then
          txc_addr_3_dly  <= '0';
        elsif set_txc_addr_3 = '1' then
          txc_addr_3_dly <= '1';
        else
          txc_addr_3_dly <= txc_addr_3_dly;
        end if;
      end if;

    end process;


    -----------------------------------------------------------------------------
    --  Generate address that will hold the End Address
    -----------------------------------------------------------------------------
    TXC_WR_ADDR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_mem_wr_addr      <= txc_min_wr_addr;
          txc_mem_wr_addr_last <= txc_wr_addr3;
          txc_mem_wr_addr_0    <= txc_wr_addr5;
          txc_mem_wr_addr_1    <= txc_wr_addr6;
        else
          if set_txc_addr_3 = '1' then
            --  increment the address for the next packet
            --  use the delayed signal to increment after the current address
            --  can be written
            if txc_mem_wr_addr = txc_max_wr_addr then
              --  if the max address is reached, loop to address 0x4
              txc_mem_wr_addr      <= txc_mem_wr_addr_0;
              txc_mem_wr_addr_last <= txc_wr_addr3;
              txc_mem_wr_addr_0    <= txc_mem_wr_addr_1;  --plus1
              txc_mem_wr_addr_1    <= txc_wr_addr6;       --plus2
            else
              --  otherwise just increment it
              txc_mem_wr_addr      <= txc_mem_wr_addr_0;
              txc_mem_wr_addr_last <= txc_mem_wr_addr;
              txc_mem_wr_addr_0    <= txc_mem_wr_addr_1;
              txc_mem_wr_addr_1    <= std_logic_vector(unsigned(txc_mem_wr_addr_1) + 1);
            end if;
          else -- Hold the current address until something changes
            txc_mem_wr_addr      <= txc_mem_wr_addr;
            txc_mem_wr_addr_last <= txc_mem_wr_addr_last;
            txc_mem_wr_addr_0    <= txc_mem_wr_addr_0;
            txc_mem_wr_addr_1    <= txc_mem_wr_addr_1;
          end if;
        end if;
      end if;
    end process;




    -----------------------------------------------------------------------------
    -- Delay the enable to align with the Memory address
    -----------------------------------------------------------------------------
    TXC_ADDR_0_DELAY : process (AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        txc_addr_0_dly1 <= set_txc_addr_0;
        txc_addr_0_dly2 <= txc_addr_0_dly1;
      end if;

    end process;


    -----------------------------------------------------------------------------
    --  Generate address that will hold the End Address
    -----------------------------------------------------------------------------
    MEM_TXC_WR_ADDR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then

        if set_txc_addr_4_n = '1' and set_txc_we = '1' then
          -- Provide the address for the End of packet address
          Axi_Str_TxC_2_Mem_Addr_int <= txc_mem_wr_addr;
        elsif set_txc_addr_3 = '1' and set_txc_we = '1' then
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr3; --set txc wr pointer
        elsif txc_addr_2 = '1' and  (txc_we = '0' or init_bram = '1') then
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr2; --get txc rd pointer
        elsif set_txc_addr_0 = '1' and (set_txc_we = '0' or init_bram = '1') then
          --  Monitor the read pointer for a full
          --  condition in the TxD Memory
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr0;
        elsif set_txc_addr_1 = '1' then
          --  Set the TxD write pointer to
          Axi_Str_TxC_2_Mem_Addr_int <= txc_wr_addr1;
        else
          Axi_Str_TxC_2_Mem_Addr_int <= (others => '0');
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_Addr <= Axi_Str_TxC_2_Mem_Addr_int;
    txc_mem_wr_addr_plus1  <= txc_mem_wr_addr_0;
    txc_mem_wr_addr_plus2  <= txc_mem_wr_addr_1;

    -----------------------------------------------------------------------------
    --  This process remaps the strobe signal to the byte address offset minus
    --  one byte.
    -----------------------------------------------------------------------------
    END_ADDRESS_BYTE_OFFSET : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txD = '1' then
          end_addr_byte_offset <= (others => '0');
        elsif axi_str_txd_tlast_dly0 = '1' and axi_str_txd_tvalid_dly0 = '1' and
              axi_str_txd_tready_int_dly = '1' then
          case axi_str_txd_tstrb_dly0 is
            when "1111" => end_addr_byte_offset <= "11";
            when "0111" => end_addr_byte_offset <= "10";
            when "0011" => end_addr_byte_offset <= "01";
            when others => end_addr_byte_offset <= "00";
          end case;
        else
          end_addr_byte_offset <= end_addr_byte_offset;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_WR_ADDR_VALUE : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' or init_bram = '1' then
          Axi_Str_TxC_2_Mem_Din_int <= (others => '0');
        elsif set_txc_addr_4_n = '1' then
        --write the ending address of the packet to memory minus one byte
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd_2 & std_logic_vector(axi_str_txd_2_mem_addr_int) & end_addr_byte_offset;
        elsif set_txc_addr_3 = '1' then
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txc & txc_mem_wr_addr;
        else
          Axi_Str_TxC_2_Mem_Din_int <= zeroes_txd & axi_str_txd_2_mem_addr_int_plus1;
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_Din <= Axi_Str_TxC_2_Mem_Din_int;

  --  Axi_Str_TxC_2_Mem_En  <= '1';
    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if (set_txc_en = '1' and set_txc_addr_2 = '0') or
           addr_2_en = '1' or init_bram = '1' then
          Axi_Str_TxC_2_Mem_En <= '1';
        else
          Axi_Str_TxC_2_Mem_En <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXC_WR_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_we = '1' then
          Axi_Str_TxC_2_Mem_We_int(0) <= '1';
        else
          Axi_Str_TxC_2_Mem_We_int(0) <= '0';
        end if;
      end if;
    end process;

    Axi_Str_TxC_2_Mem_We <= Axi_Str_TxC_2_Mem_We_int;


    -----------------------------------------------------------------------------
    --  Delay set_txc_addr_2 to align with data
    -----------------------------------------------------------------------------
    TXC_ADDR2_DLY : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_2 = '1' then
          txc_addr_2  <= set_txc_addr_2;
        else
          txc_addr_2  <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay set_txc_we to align with address
    -----------------------------------------------------------------------------
    TXC_WE_DLY : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_we = '1' then
          txc_we  <= set_txc_we;
        else
          txc_we  <= '0';
        end if;
        txc_we_dly1 <= txc_we;
        txc_we_dly2 <= txc_we_dly1;

      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Delay set_txc_we to align with address
    -----------------------------------------------------------------------------
    ADDR2_MEM_EN : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if set_txc_addr_2 = '1' and  set_txc_en = '1' then
          addr_2_en  <= set_txc_en;
        else
          addr_2_en  <= '0';
        end if;
        addr_2_en_dly1 <= addr_2_en;
        addr_2_en_dly2 <= addr_2_en_dly1;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Get the read pointer to check for FULL
    --  With ASYNC BRAM clock cannot read/write same address in memory at same
    --  time unless timing is met, so read until data matches
    -----------------------------------------------------------------------------
    MEM_TXC_RD_ADDR_PNTR : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          txc_rd_addr2_pntr_1 <= (others => '0');
          txc_rd_addr2_pntr   <= txc_min_wr_addr;
          compare_addr2_cmplt <= '0';
          compare_addr2_cmplt_dly <= '0';
        else

          if set_txc_addr_2 = '1' and addr_2_en_dly2 = '1' and txc_we_dly2 = '0' then
            txc_rd_addr2_pntr_1 <= Axi_Str_TxC_2_Mem_Dout(c_TxC_addrb_width -1 downto 0);

            if Axi_Str_TxC_2_Mem_Dout(c_TxC_addrb_width -1 downto 0) = txc_rd_addr2_pntr_1  and
               compare_addr2_cmplt = '0' then
              txc_rd_addr2_pntr   <= txc_rd_addr2_pntr_1;
              compare_addr2_cmplt <= '1';
            else
              txc_rd_addr2_pntr   <= txc_rd_addr2_pntr;
              compare_addr2_cmplt <= '0';
            end if;

          else
            txc_rd_addr2_pntr_1 <= txc_rd_addr2_pntr_1;
            txc_rd_addr2_pntr   <= txc_rd_addr2_pntr;
            compare_addr2_cmplt <= '0';
          end if;
          compare_addr2_cmplt_dly <= compare_addr2_cmplt;

        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Full flag indicator
    --    Does not begin comparison until 1st packet is written to memory
    -----------------------------------------------------------------------------
    TXC_FULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txc = '1' then
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
        elsif txc_mem_full = '1' and
           compare_addr2_cmplt = '1' and compare_addr2_cmplt_dly = '0' then
           --increments after it goes full, so use txc_mem_wr_addr for compare
          if txc_mem_wr_addr /= txc_rd_addr2_pntr then
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
          else
            txc_mem_full     <= txc_mem_full;
            txc_mem_not_full <= txc_mem_not_full;
          end if;
        elsif set_txc_addr_3 = '1' and set_txc_we = '1' then
          if txc_mem_wr_addr_plus1 = txc_rd_addr2_pntr then
            txc_mem_full     <= '1';
            txc_mem_not_full <= '0';
          else
            txc_mem_full     <= '0';
            txc_mem_not_full <= '1';
          end if;
        else
          txc_mem_full     <= txc_mem_full;
          txc_mem_not_full <= txc_mem_not_full;
        end if;
      end if;
    end process;

    TXC_AFULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if txc_mem_wr_addr_plus2 = txc_rd_addr2_pntr then
          txc_mem_afull     <= '1';
        else
          txc_mem_afull     <= '0';
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Throttle AXI Stream TxC
    --    Do not assert unless TxD is not in progress and the memory can
    --    accept data
    -----------------------------------------------------------------------------
    TXC_READY : process(AXI_STR_TXD_ACLK)
    begin



      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txc = '1' or clr_txc_trdy = '1' or clr_txc_trdy2 = '1' or
             set_txd_rdy = '1' or (txd_rdy = '1' and clr_txd_rdy = '0') or disable_txc_trdy = '1' or
             (AXI_STR_TXC_TLAST = '1' and AXI_STR_TXC_TVALID = '1' and axi_str_txc_tready_int = '1') or
             (compare_addr2 = '1' and axi_str_txc_tvalid_dly0 = '1' and axi_str_txc_tready_int_dly = '1') then
             --do not need compare_addr0 because will clr at TLAST
          axi_str_txc_tready_int <= '0';
        else

          if txc_addr_3_dly = '1' then
            if (txc_mem_wr_addr = txc_rd_addr2_pntr and txc_mem_full = '1') then
              axi_str_txc_tready_int <= '0';
            elsif txc_mem_wr_addr = txc_rd_addr2_pntr and
                Axi_Str_TxC_2_Mem_We_int(0) = '1' then
              axi_str_txc_tready_int <= '0';
            else
              axi_str_txc_tready_int <= axi_str_txc_tready_int;
            end if;
          elsif set_txc_trdy = '1' then
            axi_str_txc_tready_int <= '1';
          elsif set_txc_trdy2 = '1' then
          --  need to force it high after address compare and after reset
            axi_str_txc_tready_int <= '1';
          else
            axi_str_txc_tready_int <= axi_str_txc_tready_int;
          end if;
        end if;
        axi_str_txc_tready_int_dly <= axi_str_txc_tready_int;
      end if;
    end process;

    AXI_STR_TXC_TREADY <= axi_str_txc_tready_int;     --fix me  need to look at all txc control and TDX tlast

    -----------------------------------------------------------------------------
    --  Register and hold the axi_flag information and CSUM Control information
    --    axi_flag
    --      0x5 = Status control
    --      0xA = Normal control
    --      0xF = Null Control
    --    CSUM
    --      00 = No CSUM will be performed
    --      01 = Partial Checksum will be performed
    --      10 = Full checksum offloading will be performed
    -----------------------------------------------------------------------------
    CNTRL_WD0 : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          axi_flag   <= (others => '0');
        elsif set_axi_flag = '1' then
          axi_flag   <= axi_str_txc_tdata_dly0(31 downto 28);
        else
          axi_flag   <= axi_flag;
        end if;
      end if;
    end process;

    CNTRL_WD1 : process(AXI_STR_TXC_ACLK)
    begin

      if rising_edge(AXI_STR_TXC_ACLK) then
        if reset2axi_str_txc = '1' then
          csum_cntrl <= (others => '0');
        elsif set_csum_cntrl = '1' then
          csum_cntrl <= axi_str_txc_tdata_dly0 (1 downto  0);
        else
          csum_cntrl <= csum_cntrl;
        end if;
      end if;
    end process;

      ---------------------------------------------------------------------------
      --  Delay signal to load csum value in csum calculation
      ---------------------------------------------------------------------------
      CHECK_FULL_SIG : process(AXI_STR_TXC_ACLK)
      begin

        if rising_edge(AXI_STR_TXC_ACLK) then
          check_full <= set_txc_addr_4_n;
        end if;
      end process;



    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Data Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXD_CONTROL : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_tvalid_dly0 <= '0';
          axi_str_txd_tlast_dly0  <= '0';
          clr_txd_trdy            <= '0';
        else
          axi_str_txd_tvalid_dly0 <= AXI_STR_TXD_TVALID;
          axi_str_txd_tlast_dly0  <= AXI_STR_TXD_TLAST;
          if axi_str_txd_tvalid = '1' and axi_str_txd_tlast = '1' and axi_str_txd_tready_int = '1' then
            clr_txd_trdy <= '1';
          else
            clr_txd_trdy <= '0';
          end if;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    -- Register the incoming AXI Stream Data Bus and control signals
    -----------------------------------------------------------------------------
    REG_TXD_IN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_tstrb_dly0  <= AXI_STR_TXD_TSTRB;
        axi_str_txd_tdata_dly0  <= AXI_STR_TXD_TDATA;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Delay the data one more clock for BRAM
    -----------------------------------------------------------------------------
    REG_TXD_DLY0 : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
          axi_str_txd_tdata_dly1  <= axi_str_txd_tdata_dly0;
        else
          axi_str_txd_tdata_dly1  <= axi_str_txd_tdata_dly1;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  AXI Stream TX Data State Machine - combinational/combinatorial
    --    Used to provide the control to write the data to the BRAM
    --    This state machine will throttle the Transmit AXI Stream Control state
    --      machine until after the data information has been received.
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXD_CMB : process (txd_wr_cs,axi_str_txd_tvalid_dly0,
      axi_str_txd_tlast_dly0,
      axi_str_txd_tstrb_dly0,wrote_first_packet,axi_str_txd_tready_int_dly,
      txd_rd_pntr,txd_mem_full,txd_min_wr_addr,
      txd_rd_pntr_hold,txd_mem_afull,txd_rd_pntr_hold_plus3,
      compare_addr0_cmplt,
      axi_str_txd_2_mem_addr_int,txd_max_wr_addr,
      check_full,txd_max_wr_addr_minus4)
    begin

      inc_txd_wr_addr     <= '0';
      set_txd_we          <= "0000";
      set_txd_en          <= '0';
      set_first_packet    <= '0';
      set_txd_rdy         <= '0';
      clr_txd_rdy         <= '0';
      clr_full_pntr       <= '0';
      disable_txd_trdy    <= '0';
      disable_txc_trdy    <= '0';
      halt_pntr_update    <= '0';
      update_rd_pntrs     <= '0';

      case txd_wr_cs is
        when IDLE =>
          if compare_addr0_cmplt = '1' then
          --  Requirement is that the TXD and TXC interfaces use the same clock
          --    so it is OK to used the TXC signals in the TXD state machine
            set_txd_rdy <= '1';
            txd_wr_ns   <= TXD_PRM;
          else
            set_txd_rdy <= '0';
            txd_wr_ns   <= IDLE;
          end if;
        when TXD_PRM =>
--      Made change to ensure TxD Memory is never full here.
--      The memory can always accept data at the start of a transfer
          if axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
          --  delay incrementing pointer until next data
          --    Ethernet has to send 14bytes as a bare minimum, so it is
          --    guaranteed to get through this state with all of the strobes set
          --    and TLAST = '0'
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            disable_txd_trdy      <= '0';
            txd_wr_ns           <= TXD_WRT;
          else
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            disable_txd_trdy      <= '0';
            txd_wr_ns           <= TXD_PRM;
          end if;
        when  TXD_WRT =>
          if txd_mem_full = '1' and axi_str_txd_tready_int_dly = '0' then
          --memory is full when axi_str_txd_tready_int_dly = '0'
            inc_txd_wr_addr     <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_first_packet    <= '0';
            clr_txd_rdy         <= '0';
            disable_txd_trdy    <= '1';
            txd_wr_ns           <= MEM_FULL;
          elsif axi_str_txd_tvalid_dly0 = '1' and axi_str_txd_tready_int_dly = '1' then
            inc_txd_wr_addr     <= '1';
            set_txd_we          <= axi_str_txd_tstrb_dly0;
            set_txd_en          <= '1';
            if axi_str_txd_tlast_dly0 = '1' then
              if wrote_first_packet = '0' then
                set_first_packet <= '1';
              else
                set_first_packet <= '0';
              end if;

              clr_txd_rdy         <= '1';
              disable_txc_trdy    <= '1';
              disable_txd_trdy    <= '0';
              txd_wr_ns           <= WAIT_WR1;
            else
            --  received data (normal receive), so continue receiving data
              set_first_packet    <= '0';
              clr_txd_rdy         <= '0';
              disable_txd_trdy    <= '0';
              txd_wr_ns           <= TXD_WRT;
            end if;
          else
            inc_txd_wr_addr     <= '0';
            set_txd_we          <= "0000";
            set_txd_en          <= '0';
            set_first_packet    <= '0';
            clr_txd_rdy         <= '0';
            disable_txd_trdy    <= '0';
            txd_wr_ns           <= TXD_WRT;
          end if;
       when MEM_FULL =>
          --  stay here until the read pointer updates by 4 words or more.  The read side operates on bytes,
          --  the write side operates on words.
          --    The read pointer updates every 512 bytes (128 words) and at the end of a packet.
          --      The samallest packet the can be sent is 15bytes, but since the BRAM is 32 bit aligned,
          --      the read side will usually update the read pointer by a minimum of 16 bytes (4 words).  However,
          --      it can update by by less than 16 bytes (4 words).  This can occure if a packet started at read
          --      address 0x1A4 (write address 0x69), and the packet is 516 bytes in length (129 words).  Here the read pointer
          --      will update at 0x3A4 (write address 0xE9 - 128 words) then again at the end of the packet at 0x3A8
          --      (write address 0xEA).
          --        If this occures the below logic will detect it and update the read pointer, but stay in this
          --        state until the next update occurs.  The next update is guaranteed to be greater than 4 words,
          --        which will allow the full pointers to be cleared for the next packet.
          inc_txd_wr_addr     <= '0';
          set_txd_we          <= "0000";
          set_txd_en          <= '0';
          set_first_packet    <= '0';
          clr_txd_rdy         <= '0';
          if txd_rd_pntr = txd_rd_pntr_hold then
          --  stay here until an update occurs
            update_rd_pntrs  <= '0';
            disable_txd_trdy <= '1';
            clr_full_pntr    <= '0';
            txd_wr_ns        <= MEM_FULL;
          else
          --  The read pointer was updated to determine if it was updated by 4 words or more
          --    If not, update the hold pointers, but stay in this state
            if txd_rd_pntr_hold <= txd_max_wr_addr_minus4 then
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x0 - 0x1FB
              if txd_rd_pntr > txd_rd_pntr_hold_plus3 then
              -- an update of 4 words or greater occured so exit this state
                update_rd_pntrs  <= '0';
                disable_txd_trdy <= '0';
                clr_full_pntr    <= '1';
                txd_wr_ns        <= TXD_WRT;
              else
              --  the update was less than 4 words
              --    (txd_rd_pntr <= txd_rd_pntr_hold_plus3)
                if txd_rd_pntr < txd_rd_pntr_hold then
                --  the read pointer wrapped, so exit because the update was > 4 words
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              end if;
            else
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x1FC- 0x1FF
              if txd_rd_pntr_hold_plus3 = txd_max_wr_addr then
              --  txd_rd_pntr = 0x1FC for 2048 byte memory, so txd_rd_pntr_hold_plus3 = max memory size
                if (txd_rd_pntr <= txd_rd_pntr_hold) then
                --  the update was >= 4 words so exit
                --    for a 2048 memory, txd_rd_pntr_hold = 0x1FC
                --      if txd_rd_pntr is between 0x0 and 0x1FB then an update of 4 or more words occurred
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              else
              --  txd_rd_pntr = 0x1FD, 0x1FE, or 0x1FF for 2048 byte memory,
              --  so the minimum txd_rd_pntr_hold_plus3 can be is 0, 1, or 2
                if (txd_rd_pntr > txd_rd_pntr_hold_plus3) and (txd_rd_pntr < txd_rd_pntr_hold) then
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr has to be tween 0x1 and 0x1FC to exit this state
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr has to be tween 0x2 and 0x1FD to exit this state
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr has to be tween 0x3 and 0x1FE to exit this state
                  update_rd_pntrs  <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  txd_wr_ns        <= TXD_WRT;
                else
                --  txd_rd_pntr did not update by 4 or more words, so update hold poointers and stay in this state
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited BUT
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr was only updated 1-3 words to 0x1FE, 0x1FF, or 0x0, so stay here
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr was only updated 1-3 words to 0x1FF, 0x0, or 0x1, so stay here
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr was only updated 1-3 words to 0x0, 0x1, or 0x2, so stay here
                  update_rd_pntrs  <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= MEM_FULL;
                end if;
              end if;
            end if;
          end if;

        when WAIT_WR1 =>
          disable_txc_trdy  <= '1';
          disable_txd_trdy  <= '0';

          if check_full = '1' then
            txd_wr_ns         <= WAIT_WR2;
          else
            txd_wr_ns         <= WAIT_WR1;
          end if;
        when WAIT_WR2 =>
          if txd_mem_full = '1' or txd_mem_afull = '1' then
            disable_txc_trdy  <= '1';
            disable_txd_trdy  <= '1';
            txd_wr_ns         <= CLR_FULL;
          else
            if wrote_first_packet = '0' then
              set_first_packet <= '1';
            else
              set_first_packet <= '0';
            end if;

            disable_txc_trdy  <= '0';
            disable_txd_trdy  <= '0';
            txd_wr_ns         <= IDLE;
          end if;

        when CLR_FULL =>
          --  stay here until the read pointer updates by 4 words or more.  The read side operates on bytes,
          --  the write side operates on words.
          --    The read pointer updates every 512 bytes (128 words) and at the end of a packet.
          --      The samallest packet the can be sent is 15bytes, but since the BRAM is 32 bit aligned,
          --      the read side will usually update the read pointer by a minimum of 16 bytes (4 words).  However,
          --      it can update by by less than 16 bytes (4 words).  This can occure if a packet started at read
          --      address 0x1A4 (write address 0x69), and the packet is 516 bytes in length (129 words).  Here the read pointer
          --      will update at 0x3A4 (write address 0xE9 - 128 words) then again at the end of the packet at 0x3A8
          --      (write address 0xEA).
          --        If this occures the below logic will detect it and update the read pointer, but stay in this
          --        state until the next update occurs.  The next update is guaranteed to be greater than 4 words,
          --        which will allow the full pointers to be cleared for the next packet.
          inc_txd_wr_addr     <= '0';
          set_txd_we          <= "0000";
          set_txd_en          <= '0';
          set_first_packet    <= '0';
          clr_txd_rdy         <= '0';
          if txd_rd_pntr = txd_rd_pntr_hold then
          --  stay here until an update occurs
            update_rd_pntrs  <= '0';
            halt_pntr_update <= '1';
            disable_txc_trdy <= '1';
            disable_txd_trdy <= '1';
            clr_full_pntr    <= '0';
            txd_wr_ns        <= CLR_FULL;
          else
          --  The read pointer was updated to determine if it was updated by 4 words or more
          --    If not, update the hold pointers, but stay in this state
            if txd_rd_pntr_hold <= txd_max_wr_addr_minus4 then
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x0 - 0x1FB
              if txd_rd_pntr > txd_rd_pntr_hold_plus3 then
              -- an update of 4 words or greater occured so exit this state
                if wrote_first_packet = '0' then
                  set_first_packet <= '1';
                else
                  set_first_packet <= '0';
                end if;
                update_rd_pntrs  <= '0';
                halt_pntr_update <= '0';
                disable_txd_trdy <= '0';
                clr_full_pntr    <= '1';
                clr_txd_rdy      <= '0';
                txd_wr_ns        <= WAIT_COMPARE_CMPLT;
              else
              --  the update was less than 4 words
              --    (txd_rd_pntr <= txd_rd_pntr_hold_plus3)
                if txd_rd_pntr < txd_rd_pntr_hold then
                --  the read pointer wrapped, so exit because the update was > 4 words
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  halt_pntr_update <= '1';
                  disable_txc_trdy <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= CLR_FULL;
                end if;
              end if;
            else
            --  for 2048 mem this covers from txd_rd_pntr_hold = 0x1FC- 0x1FF
              if txd_rd_pntr_hold_plus3 = txd_max_wr_addr then
              --  txd_rd_pntr = 0x1FC for 2048 byte memory, so txd_rd_pntr_hold_plus3 = max memory size
                if (txd_rd_pntr <= txd_rd_pntr_hold) then
                --  the update was >= 4 words so exit
                --    for a 2048 memory, txd_rd_pntr_hold = 0x1FC
                --      if txd_rd_pntr is between 0x0 and 0x1FB then an update of 4 or more words occurred
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  the update was less than 4 words, so update the read hold pointers and stay here until the next update
                --    txd_rd_pntr >= txd_rd_pntr_hold
                  update_rd_pntrs  <= '1';
                  halt_pntr_update <= '1';
                  disable_txc_trdy <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= CLR_FULL;
                end if;
              else
              --  txd_rd_pntr = 0x1FD, 0x1FE, or 0x1FF for 2048 byte memory,
              --  so the minimum txd_rd_pntr_hold_plus3 can be is 0, 1, or 2
                if (txd_rd_pntr > txd_rd_pntr_hold_plus3) and (txd_rd_pntr < txd_rd_pntr_hold) then
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr has to be tween 0x1 and 0x1FC to exit this state
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr has to be tween 0x2 and 0x1FD to exit this state
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr has to be tween 0x3 and 0x1FE to exit this state
                  if wrote_first_packet = '0' then
                    set_first_packet <= '1';
                  else
                    set_first_packet <= '0';
                  end if;
                  update_rd_pntrs  <= '0';
                  halt_pntr_update <= '0';
                  disable_txd_trdy <= '0';
                  clr_full_pntr    <= '1';
                  clr_txd_rdy      <= '0';
                  txd_wr_ns        <= WAIT_COMPARE_CMPLT;
                else
                --  txd_rd_pntr did not update by 4 or more words, so update hold poointers and stay in this state
                --  txd_rd_pntr_hold will be either 0x1FD, 0x1FE, or 0x1FF for a 2048 byte memory
                --    if txd_rd_pntr >  txd_rd_pntr_hold and  txd_rd_pntr <  txd_rd_pntr_hold
                --      then the update was >= 4 words and the state can be exited BUT
                --          if  txd_rd_pntr_hold = 0x1FD then  txd_rd_pntr_hold_plus3 = 0
                --            txd_rd_pntr was only updated 1-3 words to 0x1FE, 0x1FF, or 0x0, so stay here
                --          if  txd_rd_pntr_hold = 0x1FE then  txd_rd_pntr_hold_plus3 = 1
                --            txd_rd_pntr was only updated 1-3 words to 0x1FF, 0x0, or 0x1, so stay here
                --          if  txd_rd_pntr_hold = 0x1FF then  txd_rd_pntr_hold_plus3 = 2
                --            txd_rd_pntr was only updated 1-3 words to 0x0, 0x1, or 0x2, so stay here
                  update_rd_pntrs  <= '1';
                  halt_pntr_update <= '1';
                  disable_txc_trdy <= '1';
                  disable_txd_trdy <= '1';
                  clr_full_pntr    <= '0';
                  txd_wr_ns        <= CLR_FULL;
                end if;
              end if;
            end if;
          end if;

        when WAIT_COMPARE_CMPLT =>
          txd_wr_ns        <= IDLE;
        when others =>
          txd_wr_ns <= IDLE;
      end case;
    end process;

    -----------------------------------------------------------------------------
    -- AXI Stream TX Control State Machine Sequencer
    -----------------------------------------------------------------------------
    FSM_AXISTRM_TXD_SEQ : process (AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_wr_cs <= IDLE;
        else
          txd_wr_cs <= txd_wr_ns;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    -- Indicator when performing a write to TxD Memory
    --  clear on axi_str_txd_tlast_dly0 = '1'
    -----------------------------------------------------------------------------
    TXD_RDY_INDICATOR : process (AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rdy <= '0';
        else
          if clr_txd_rdy = '1' then
            txd_rdy <= '0';
          elsif set_txd_rdy = '1' then
            txd_rdy <= '1';
          else
            txd_rdy <= txd_rdy;
          end if;
        end if;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Filter to indicate first packet was written
    --    Needed for full flag
    -----------------------------------------------------------------------------
    FIRST_PACKET_WROTE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          wrote_first_packet <= '0';
        elsif set_first_packet = '1' then
          wrote_first_packet <= '1';
        else
          wrote_first_packet <= wrote_first_packet;
        end if;
      end if;
    end process;


    axi_str_txd_2_mem_addr_int_plus1 <= std_logic_vector(axi_str_txd_2_mem_addr_int + 1);
    axi_str_txd_2_mem_addr_int_plus2 <= std_logic_vector(axi_str_txd_2_mem_addr_int + 2);
    axi_str_txd_2_mem_addr_int_plus3 <= std_logic_vector(axi_str_txd_2_mem_addr_int + 3);
    axi_str_txd_2_mem_addr_int_plus4 <= std_logic_vector(axi_str_txd_2_mem_addr_int + 4);


    ---------------------------------------------------------------------------
    --  Register to help fmax
    --  With ASYNC BRAM clock cannot read/write same address in memory at same
    --  time unless timing is met, so read until data matches
    ---------------------------------------------------------------------------
    RD_PNTR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rd_pntr_1 <= (others => '0');
          txd_rd_pntr   <= (others => '0');
          compare_addr0_cmplt <= '0';
        else
          if set_txc_addr_0 = '1' and txc_addr_0_dly2 = '1' and
             txc_we_dly2 = '0'  then
          --  txc_addr_0_dly2 is when data is first avaliable from memory

          --  use set_txc_addr_0 to disable compare_addr0_cmplt once pointers update
          --  once state machine advances, set_txc_addr_0 will go low so use it to disable any more
          --  any more data from memory
            txd_rd_pntr_1      <= Axi_Str_TxC_2_Mem_Dout(c_TxD_addrb_width -1 downto 0);

            if Axi_Str_TxC_2_Mem_Dout(c_TxD_addrb_width -1 downto 0) = txd_rd_pntr_1 and
              compare_addr0_cmplt = '0' then
              txd_rd_pntr         <= txd_rd_pntr_1;
              if enable_compare_addr0_cmplt = '1' then
                compare_addr0_cmplt <= '1';
              else
                compare_addr0_cmplt <= '0';
              end if;
            else
              txd_rd_pntr         <= txd_rd_pntr;
              compare_addr0_cmplt <= '0';
            end if;
          else
            txd_rd_pntr_1      <= txd_rd_pntr_1;
            txd_rd_pntr        <= txd_rd_pntr;
            compare_addr0_cmplt<= '0';
          end if;
        end if;
      end if;
    end process;


    ---------------------------------------------------------------------------
    --  Update the read pointer locations until the memory goes FULL
    --    Then use the stored values to compare against real time read pointer
    --    and throttle appropriately
    ---------------------------------------------------------------------------
    RD_PNTRS : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          txd_rd_pntr_hold_plus3 <= txc_rd_addr3;
          txd_rd_pntr_hold       <= txc_rd_addr0;
        else
          if (txd_mem_full = '0' and txc_addr_0_dly2 = '1' and halt_pntr_update = '0') or update_rd_pntrs = '1'then -- wait on this as it might not be needed  or update_hold_pntrs = '1' then --and
          --  halt_pntr_update is for the special case when memory is almost full/full and
          --  the Txd FSM needs to wait for a few reads before the next packet starts
          --  The TxD FSM will assert it HIGH to prevent the poiners from being updated
            txd_rd_pntr_hold_plus3 <= std_logic_vector(unsigned(txd_rd_pntr) +3);
            txd_rd_pntr_hold       <= txd_rd_pntr;
          else
            txd_rd_pntr_hold_plus3 <= txd_rd_pntr_hold_plus3;
            txd_rd_pntr_hold       <= txd_rd_pntr_hold;
          end if;
        end if;
      end if;
    end process;


    -----------------------------------------------------------------------------
    --  Full flag indicator
    --    Does not begin comparison until 1st packet is written to memory
    -----------------------------------------------------------------------------
    TXD_FULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
            txd_mem_full     <= '0';
            txd_mem_not_full <= '1';
        else
            if (axi_str_txd_2_mem_addr_int_plus3 = txd_rd_pntr and
              (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) then
              txd_mem_full     <= '1';
              txd_mem_not_full <= '0';
            else
              txd_mem_full     <= txd_mem_full;
              txd_mem_not_full <= txd_mem_not_full;
            end if;
        end if;
      end if;
    end process;

    TXD_AFULL_FLAG : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_full_pntr = '1' then
            txd_mem_afull     <= '0';
        else

          if (axi_str_txd_2_mem_addr_int_plus4 = txd_rd_pntr and
              (inc_txd_wr_addr = '1'  or inc_txd_addr_one = '1')) then
            txd_mem_afull     <= '1';
          else
            txd_mem_afull     <= txd_mem_afull;
          end if;
        end if;
      end if;
    end process;

    DELAY_TXD_TREADY_DISABLE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        disable_txd_trdy_dly <= disable_txd_trdy;
      end if;
    end process;

    DELAY_TREADY_DISABLE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        disable_txc_trdy_dly <= disable_txc_trdy;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  TxD Ready
    --    Only assert when FIFO is not full and TxC is not in process
    -----------------------------------------------------------------------------
    TXD_READY : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_tready_int_dly <= axi_str_txd_tready_int;
        if (AXI_STR_TXD_TLAST = '1' and AXI_STR_TXD_TVALID = '1' and axi_str_txd_tready_int = '1') or
           (clr_txd_trdy = '1' and disable_txd_trdy_dly = '0') or
           disable_txd_trdy = '1' then
          axi_str_txd_tready_int <= '0';
        elsif set_txd_rdy = '1' or (txd_rdy = '1' and clr_txd_rdy = '0') then
            if (axi_str_txd_2_mem_addr_int_plus3 = txd_rd_pntr and
               inc_txd_wr_addr = '1') or
               (clr_full_pntr = '0' and txd_mem_full = '1') then
            --  txd_rd_pntr is where the the current read is occuring, so
            --    to account for register pipelines, this needs to stop at
            --    3 counts before the current write address
              axi_str_txd_tready_int <= '0';
            else
              axi_str_txd_tready_int <= '1';
            end if;
        else
          axi_str_txd_tready_int <= '0';
        end if;
      end if;
    end process;

    AXI_STR_TXD_TREADY     <= axi_str_txd_tready_int;    --fix me  need to look at all txd control and TXC tlast

    -----------------------------------------------------------------------------
    --  Address to AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_WR_ADDR : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' then
          axi_str_txd_2_mem_addr_int <= (others => '0');
        elsif (inc_txd_wr_addr = '1' or inc_txd_addr_one = '1') then
        --  the address ready for the next transaction
          axi_str_txd_2_mem_addr_int <= axi_str_txd_2_mem_addr_int + 1;
        else
          axi_str_txd_2_mem_addr_int <= axi_str_txd_2_mem_addr_int;
        end if;
      end if;
    end process;

    ---------------------------------------------------------------------------
    --  Force and update the BRAM with the axi_str_txd_2_mem_addr_int
    --  every ~128 writes (~512 bytes)
    ---------------------------------------------------------------------------
    BRAM_UPDATE : process(AXI_STR_TXD_ACLK)
    begin

      if rising_edge(AXI_STR_TXD_ACLK) then
        if reset2axi_str_txd = '1' or clr_txd_rdy = '1' then
          update_bram_cnt     <= (others => '0');
        else
          if update_bram_cnt(7) = '1' and inc_txd_wr_addr = '1' then
            update_bram_cnt <= std_logic_vector(unsigned('0' & update_bram_cnt(6 downto 0)) + 1);
          elsif inc_txd_wr_addr = '1' then
            update_bram_cnt <= std_logic_vector(unsigned(update_bram_cnt) + 1);
          else
            update_bram_cnt <= update_bram_cnt;
          end if;
        end if;
      end if;
    end process;


    axi_str_txd_2_mem_addr               <= std_logic_vector(axi_str_txd_2_mem_addr_int);


    Axi_Str_TxD_2_Mem_Din(35)           <= axi_str_txd_2_mem_we_int(3);
    Axi_Str_TxD_2_Mem_Din(26)           <= axi_str_txd_2_mem_we_int(2);
    Axi_Str_TxD_2_Mem_Din(17)           <= axi_str_txd_2_mem_we_int(1);
    Axi_Str_TxD_2_Mem_Din(8)            <= axi_str_txd_2_mem_we_int(0);

    Axi_Str_TxD_2_Mem_Din(34 downto 27) <= axi_str_txd_tdata_dly1(31 downto 24);
    Axi_Str_TxD_2_Mem_Din(25 downto 18) <= axi_str_txd_tdata_dly1(23 downto 16);
    Axi_Str_TxD_2_Mem_Din(16 downto  9) <= axi_str_txd_tdata_dly1(15 downto  8);
    Axi_Str_TxD_2_Mem_Din(7  downto  0) <= axi_str_txd_tdata_dly1( 7 downto  0);

    -----------------------------------------------------------------------------
    --  Write Parity bits to the AXI Stream Data Memory
    --    The parity bit always should be the AXI_STR_TXD_TSTRB bits delayed
    -----------------------------------------------------------------------------
    MEM_TXD_PARITY : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        axi_str_txd_2_mem_we_int <= set_txd_we;
      end if;
    end process;

    -----------------------------------------------------------------------------
    --  Write Enable bits to the AXI Stream Data Memory
    --    All of the write enables bits should be forced HIGH any time a write to
    --    memory is being performed.  This will allow the parity bits to be
    --    cleared which in turn prevents too much data being read on the Txd
    --    client interface.
    -----------------------------------------------------------------------------
    MEM_TXD_WR_EN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        case set_txd_we is
          when "0000" => Axi_Str_TxD_2_Mem_We <= "0000";
          when others => Axi_Str_TxD_2_Mem_We <= "1111";
        end case;
      end if;
    end process;

--    Axi_Str_TxD_2_Mem_We <= axi_str_txd_2_mem_we_int;

    -----------------------------------------------------------------------------
    --  Enable bit to the AXI Stream Data Memory
    -----------------------------------------------------------------------------
    MEM_TXD_EN : process(AXI_STR_TXD_ACLK)
    begin
      if rising_edge(AXI_STR_TXD_ACLK) then
        if set_txd_en = '1' then
          axi_str_txd_2_mem_en_int <= '1';
        else
          axi_str_txd_2_mem_en_int <= '0';
        end if;
      end if;
    end process;

    Axi_Str_TxD_2_Mem_En <= axi_str_txd_2_mem_en_int;

-------------------------------------------------------------------------------
--  End Basic Design
-------------------------------------------------------------------------------

end rtl;


-------------------------------------------------------------------------------
-- tx_emac_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename: tx_emac_if.vhd
-- Version: v1.00a
-- Description: top level of embedded ip Ethernet MAC interface
--
-- VHDL-Standard: VHDL'93
-------------------------------------------------------------------------------
-- Structure: This section shows the hierarchical structure of axi_ethernet.
--
-- axi_ethernet.vhd
-- axi_ethernt_soft_temac_wrap.vhd
-- axi_lite_ipif.vhd
-- embedded_top.vhd
-- tx_if.vhd
-- tx_axistream_if.vhd
-- tx_mem_if
-- -> tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author: MW
--
-- MW 07/01/10
-- ^^^^^^
-- - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
-- active low signals: "*_n"
-- clock signals: "clk", "clk_div#", "clk_#x"
-- reset signals: "rst", "rst_n"
-- generics: "C_*"
-- user defined types: "*_TYPE"
-- state machine next state: "*_ns"
-- state machine current state: "*_cs"
-- combinatorial signals: "*_com"
-- pipelined or register delay signals: "*_d#"
-- counter signals: "*cnt*"
-- clock enable signals: "*_ce"
-- internal version of output port "*_i"
-- device pins: "*_pin"
-- ports: - Names begin with Uppercase
-- processes: "*_PROCESS"
-- component instantiations: "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tx_if_pack.all;


-------------------------------------------------------------------------------
-- Entity Section
-------------------------------------------------------------------------------

entity tx_emac_if is
  generic (
    C_FAMILY            : string                   := "virtex6";
    C_HALFDUP           : integer range 0 to 1     := 0;
    C_TXMEM             : integer                  := 4096;
    C_TXCSUM            : integer range 0 to 2     := 0;
    C_ENABLE_1588       : integer                  := 0;

-- Read Port - AXI Stream TxData
    c_TxD_write_width_a : integer range 0 to 18    := 9;
    c_TxD_read_width_a  : integer range 0 to 18    := 9;
    c_TxD_write_depth_a : integer range 0 to 32768 := 4096;
    c_TxD_read_depth_a  : integer range 0 to 32768 := 4096;
    c_TxD_addra_width   : integer range 0 to 15    := 10;
    c_TxD_wea_width     : integer range 0 to 2     := 2;

-- Read Port - AXI Stream TxControl
    c_TxC_write_width_a : integer range 36 to 36   := 36;
    c_TxC_read_width_a  : integer range 36 to 36   := 36;
    c_TxC_write_depth_a : integer range 0 to 1024  := 1024;
    c_TxC_read_depth_a  : integer range 0 to 1024  := 1024;
    c_TxC_addra_width   : integer range 0 to 10    := 10;
    c_TxC_wea_width     : integer range 0 to 1     := 1;

    c_TxD_addrb_width   : integer range 0 to 13    := 10;

    C_CLIENT_WIDTH      : integer                  := 8
    );
  port (
--Transmit Memory Read Interface
-- ** WARNING ** WARNING ** WARNING **
--  For MII,GMII, RGMI, 1000Base-X and pcs/pma SGMII this is an accurate indicator
--  However for V6 Hard SGMII it is always tied to '0' for all speeds
    tx_client_10_100         : in  std_logic; --  Tx Client CE Toggles Indicator

-- Read Port - AXI Stream TxData
    reset2tx_client          : in  std_logic; --  reset
    Tx_Client_TxD_2_Mem_Din  : out std_logic_vector (c_TxD_write_width_a-1 downto 0); --  Tx AXI-Stream Data to Memory Wr Din
    Tx_Client_TxD_2_Mem_Addr : out std_logic_vector (c_TxD_addra_width-1 downto 0  ); --  Tx AXI-Stream Data to Memory Wr Addr
    Tx_Client_TxD_2_Mem_En   : out std_logic; --  Tx AXI-Stream Data to Memory Enable
    Tx_Client_TxD_2_Mem_We   : out std_logic_vector (c_TxD_wea_width-1 downto 0    ); --  Tx AXI-Stream Data to Memory Wr En
    Tx_Client_TxD_2_Mem_Dout : in  std_logic_vector (c_TxD_read_width_a-1 downto 0 ); --  Tx AXI-Stream Data to Memory Not Used

-- Read Port - AXI Stream TxControl
    reset2axi_str_txd        : in  std_logic; --  reset
    Tx_Client_TxC_2_Mem_Din  : out std_logic_vector (c_TxC_write_width_a-1 downto 0); --  Tx AXI-Stream Control to Memory Wr Din
    Tx_Client_TxC_2_Mem_Addr : out std_logic_vector (c_TxC_addra_width-1 downto 0  ); --  Tx AXI-Stream Control to Memory Wr Addr
    Tx_Client_TxC_2_Mem_En   : out std_logic; --  Tx AXI-Stream Control to Memory Enable
    Tx_Client_TxC_2_Mem_We   : out std_logic_vector (c_TxC_wea_width-1 downto 0    ); --  Tx AXI-Stream Control to Memory Wr En
    Tx_Client_TxC_2_Mem_Dout : in  std_logic_vector (c_TxC_read_width_a-1 downto 0 ); --  Tx AXI-Stream Control to Memory Full Flag

--  Tx AXI-S Interface
    tx_axi_clk               : in  std_logic; --  Tx AXI-Stream clock in
    tx_reset_out             : in  std_logic; --  take to reset combiner
    tx_axis_mac_tdata        : out std_logic_vector (C_CLIENT_WIDTH - 1 downto 0   ); --  Tx AXI-Stream data
    tx_axis_mac_tvalid       : out std_logic; --  Tx AXI-Stream valid
    tx_axis_mac_tlast        : out std_logic; --  Tx AXI-Stream last
    tx_axis_mac_tuser        : out std_logic; -- this is always driven low since an underflow cannot occur
    tx_axis_mac_tready       : in  std_logic; --  Tx AXI-Stream ready in from TEMAC
    tx_collision             : in  std_logic; --  collision not used
    tx_retransmit            : in  std_logic; -- retransmit not used


    tx_cmplt                 : out std_logic; -- transmit is complete indicator

    tx_init_in_prog_cross    : in  std_logic        --  Tx is Initializing after a reset
    );

end tx_emac_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of tx_emac_if is

    type TXC_RD_FSM_TYPE is (
    GET_TXC_WR_PNTR,
    GET_END_PNTR,
    SET_TXCRD_PNTR,
    GET_TXDWR_PNTR,
    SET_TXDRD_PNTR,
    WAIT_TXD_DONE,
    GET_ADDR3,
    WAIT_ADDR3_PNTR);

    signal txc_rd_cs, txc_rd_ns : TXC_RD_FSM_TYPE;

    type TXD_RD_FSM_TYPE is (
    IDLE,
    GET_1588_CMD1,
    GET_1588_CMD2,
    GET_1588_CMD3,
    GET_1588_CMD4,
    GET_1588_CMD5,
    GET_1588_CMD6,
    GET_1588_CMD7,
    GET_1588_CMD8,
    GET_B1,
    GET_B2,
    GET_B3,
    GET_B4,
    WAIT_TRDY2,
    WAIT_TRDY3,
    PRM_DATA,
    CHECK_DONE,
    WAIT_LAST);

    signal txd_rd_cs, txd_rd_ns : TXD_RD_FSM_TYPE;

    signal enable_1588_val     : std_logic_vector(2 downto 0) := (others => '0'); 
    signal enabled_1588        : std_logic;
    signal set_txc_addr0       : std_logic;
    signal set_txc_addr1       : std_logic;
    signal set_txc_addr2       : std_logic;
    signal set_txc_addr3       : std_logic;
    signal set_txc_addr3_d1    : std_logic;
    signal txc_addr3_en        : std_logic;
    signal set_txc_addr4_n     : std_logic;
    signal set_txc_wr          : std_logic;
    signal set_txc_en          : std_logic;
    signal txc_wr_pntr_en      : std_logic;
    signal set_start_txd_fsm   : std_logic;
    signal start_txd_fsm       : std_logic;
    signal inc_txc_rd_addr     : std_logic;
    signal first_rd            : std_logic;
    signal txc_wr_pntr_1       : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_wr_pntr_2       : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_wr_pntr         : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal compare_addr3_cmplt : std_logic;

    signal Tx_Client_TxC_2_Mem_Addr_int : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_mem_rd_addr              : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr_cmp              : std_logic_vector(c_TxC_addra_width -1 downto 0);

    signal end_addr                    : std_logic_vector(c_TxD_addra_width -1 downto 0);
    signal txc_rd_end                  : std_logic;
    signal txc_rd_end_dly1             : std_logic;
    signal Tx_Client_TxC_2_Mem_En_int  : std_logic;
    signal Tx_Client_TxC_2_Mem_We_int  : std_logic_vector(c_TxC_wea_width-1 downto 0);
    signal Tx_Client_TxC_2_Mem_Din_int : std_logic_vector(c_TxC_write_width_a -1 downto 0);

    signal set_txd_vld            : std_logic;
    signal set_txd_vld_1          : std_logic;
    signal set_txd_vld_2          : std_logic;
    signal clr_txd_vld            : std_logic;
    signal set_txd_en             : std_logic;
    signal inc_txd_rd_addr        : std_logic;
    signal txd_rd_addr            : std_logic_vector(c_TxD_addra_width -1 downto 0);
    signal txd_rd_addr_1_0        : std_logic_vector(1 downto 0);
    signal txd_rd_addr_aligned    : std_logic_vector(c_TxD_addra_width -1 downto 0);
    signal txd_wr_pntr_en         : std_logic;

    signal align_start_addr           : std_logic;
    signal set_txd_done               : std_logic;
    signal Tx_Client_TxD_2_Mem_En_int : std_logic;
    signal txd                        : std_logic_vector(C_CLIENT_WIDTH-1 downto 0);
    signal txd_vld                    : std_logic;

    signal txc_min_rd_addr : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_max_rd_addr : std_logic_vector(c_TxC_addra_width -1 downto 0);

    signal txc_rd_addr0 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr1 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr2 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr3 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr5 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr6 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr7 : std_logic_vector(c_TxC_addra_width -1 downto 0);

    signal txc_mem_rd_addr_0 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_mem_rd_addr_1 : std_logic_vector(c_TxC_addra_width -1 downto 0);

    signal txd_1 : std_logic_vector(C_CLIENT_WIDTH-1 downto 0);
    signal txd_2 : std_logic_vector(C_CLIENT_WIDTH-1 downto 0);
    signal txd_3 : std_logic_vector(C_CLIENT_WIDTH-1 downto 0);

    constant zeroes_txc : std_logic_vector(c_TxC_read_width_a -1 downto c_TxC_addra_width)    := (others => '0');
    constant zeroes_txd : std_logic_vector(c_TxC_read_width_a -1 downto c_TxD_addra_width -2) := (others => '0');

    signal txcl_init_in_prog_dly1 : std_logic;
    signal txcl_init_in_prog_dly2 : std_logic;
    signal txcl_init_in_prog_dly3 : std_logic;
    signal txcl_init_in_prog_dly4 : std_logic;

    signal update_bram_cnt : unsigned(9 downto 0);

    signal tx_axis_mac_tready_dly : std_logic;
    signal mux_b3                 : std_logic;

    signal tx_axis_mac_tlast_int : std_logic;

    signal set_byte_en      : std_logic;
    signal set_byte_en_pipe : std_logic_vector(1 downto 0);
    signal set_first_bytes  : std_logic;
    signal first_bytes      : std_logic;

    signal phy_mode_enable : std_logic;

begin

    tx_axis_mac_tuser <= '0';

    Tx_Client_TxD_2_Mem_Din <= (others => '0');

    phy_mode_enable <= tx_client_10_100;

    enable_1588_val <= std_logic_vector(to_unsigned(C_ENABLE_1588, enable_1588_val'length));
    enabled_1588 <= '1' when ((enable_1588_val(1) = '1' and enable_1588_val(0) = '0') or (enable_1588_val(1) = '0' and enable_1588_val(0) = '1')) 
                    else '0';

-----------------------------------------------------------------------------
--  Create the full and empty comparison values for the S6 and V6 since
--  1 S6 BRAM = 1/2 V6 BRAM
-----------------------------------------------------------------------------
    GEN_TXC_MIN_MAX_RD_FLAG : for i in (c_TxC_addra_width - 1) downto 0 generate
        txc_min_rd_addr(i) <= '1' when (i = 2)                   else '0';
        txc_max_rd_addr(i) <= '0' when (i = 0 or i = 1)          else '1';
        txc_rd_addr0(i)    <= '0';
        txc_rd_addr1(i)    <= '1' when (i = 0)                   else '0';
        txc_rd_addr2(i)    <= '1' when (i = 1)                   else '0';
        txc_rd_addr3(i)    <= '1' when (i = 0 or i = 1)          else '0';
        txc_rd_addr5(i)    <= '1' when (i = 0 or i = 2)          else '0';
        txc_rd_addr6(i)    <= '1' when (i = 1 or i = 2)          else '0';
        txc_rd_addr7(i)    <= '1' when (i = 0 or i = 1 or i = 2) else '0';

    end generate GEN_TXC_MIN_MAX_RD_FLAG;

-----------------------------------------------------------------------------
--  Transmit Client TX Control State Machine Combinatorial Logic
-----------------------------------------------------------------------------
    FSM_TXCLIENT_TXC_CMB : process (txc_rd_cs,tx_axis_mac_tready,
      clr_txd_vld,txc_rd_addr_cmp,
      txcl_init_in_prog_dly4,compare_addr3_cmplt,txc_wr_pntr,
      update_bram_cnt)
    begin
        set_txc_addr0     <= '0';
        set_txc_addr1     <= '0';
        set_txc_addr2     <= '0';
        set_txc_addr3     <= '0';
        set_txc_addr4_n   <= '0';
        set_txc_wr        <= '0';
        set_txc_en        <= '0';
        set_start_txd_fsm <= '0';
        inc_txc_rd_addr   <= '0';

        case txc_rd_cs is
            when GET_TXC_WR_PNTR =>
                if txcl_init_in_prog_dly4 = '0' and compare_addr3_cmplt = '1' and txc_rd_addr_cmp /= txc_wr_pntr then
                    set_txc_addr3     <= '0';
                    set_txc_addr4_n   <= '1'; -- Read TxC Addr 0x4 - 0xn
                    set_txc_en        <= '1';
                    inc_txc_rd_addr   <= '1';
                    txc_rd_ns         <= GET_END_PNTR;
                else
                    set_txc_addr3     <= '1'; -- Read TxC Addr 0x3 (TxC Empty)
                    set_txc_addr4_n   <= '0';
                    set_txc_en        <= '1';
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= GET_TXC_WR_PNTR;
                end if;
            when GET_END_PNTR    =>
                set_txc_addr2       <= '1'; -- Write TxC Addr 0x2
                set_txc_wr          <= '1';
                set_txc_en          <= '1';
                txc_rd_ns           <= SET_TXCRD_PNTR;
            when SET_TXCRD_PNTR  =>
                set_txc_addr1       <= '1'; -- Read TxC Addr 0x1
                set_txc_en          <= '1';
                txc_rd_ns           <= GET_TXDWR_PNTR;
            when GET_TXDWR_PNTR  =>
                set_txc_addr0       <= '1'; -- Write TxC Addr 0x0
                set_txc_wr          <= '1';
                set_txc_en          <= '1';
                txc_rd_ns           <= SET_TXDRD_PNTR;
            when SET_TXDRD_PNTR  =>
                set_txc_addr0       <= '0';
                set_txc_wr          <= '0';
                set_txc_en          <= '0';
                set_start_txd_fsm   <= '1';
                txc_rd_ns           <= WAIT_TXD_DONE;
            when WAIT_TXD_DONE   =>
                if tx_axis_mac_tready = '1' and clr_txd_vld = '0' then
                    if update_bram_cnt(9) = '1' then  --Update the TxC BRAM with the current rd_addr_addr
                        set_txc_addr0   <= '1'; -- Write TxC Addr 0x0
                        set_txc_addr3   <= '0';
                        set_txc_wr      <= '1';
                        set_txc_en      <= '1';
                        inc_txc_rd_addr <= '0';
                        txc_rd_ns       <= WAIT_TXD_DONE;
                    else
                        set_txc_addr0   <= '0'; -- Write TxC Addr 0x0
                        set_txc_addr3   <= '0';
                        set_txc_wr      <= '0';
                        set_txc_en      <= '0';
                        inc_txc_rd_addr <= '0';
                        txc_rd_ns       <= WAIT_TXD_DONE;
                    end if;
                elsif tx_axis_mac_tready = '1' and clr_txd_vld = '1' then
                    set_txc_addr0     <= '1';
                    set_txc_addr3     <= '0';
                    set_txc_wr        <= '1';
                    set_txc_en        <= '1'; --write the last rd_rntr_addr for this packet
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= GET_ADDR3;
                else
                    set_txc_addr0     <= '0';
                    set_txc_addr3     <= '0'; --do nothing
                    set_txc_wr        <= '0';
                    set_txc_en        <= '0';
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= WAIT_TXD_DONE;
                end if;
            when GET_ADDR3       =>
                if tx_axis_mac_tready = '1' then
                    set_txc_addr0     <= '0';
                    set_txc_addr3     <= '1';
                    set_txc_wr        <= '0';
                    set_txc_en        <= '1'; --get ready for the next packet - addr0x4-0xn
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= WAIT_ADDR3_PNTR;
                else
                    set_txc_addr0     <= '0';
                    set_txc_addr3     <= '0';
                    set_txc_wr        <= '0';
                    set_txc_en        <= '0';
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= GET_ADDR3;
                end if;
            when WAIT_ADDR3_PNTR =>
                set_txc_addr0       <= '0';
                set_txc_addr3       <= '1';
                set_txc_wr          <= '0';
                set_txc_en          <= '1';
                inc_txc_rd_addr     <= '0';
                txc_rd_ns           <= GET_TXC_WR_PNTR;
            when others          =>
                txc_rd_ns           <= GET_TXC_WR_PNTR;
        end case;
    end process;

-----------------------------------------------------------------------------
--  Transmit Client TX Control State Machine Sequencer
-----------------------------------------------------------------------------
  FSM_TXCLIENT_TXC_SEQ : process (tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txc_rd_cs <= GET_TXC_WR_PNTR;
      else
        txc_rd_cs <= txc_rd_ns;
      end if;
    end if;
  end process;

---------------------------------------------------------------------------
--  Delay the indicator to ensure the memory has had enough time to update
---------------------------------------------------------------------------
  TXCL_INIT_INDICATOR_DLY : process (tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txcl_init_in_prog_dly1 <= '1';
        txcl_init_in_prog_dly2 <= '1';
        txcl_init_in_prog_dly3 <= '1';
        txcl_init_in_prog_dly4 <= '1';
      else
        txcl_init_in_prog_dly1 <= tx_init_in_prog_cross;
        txcl_init_in_prog_dly2 <= txcl_init_in_prog_dly1;
        txcl_init_in_prog_dly3 <= txcl_init_in_prog_dly2;
        txcl_init_in_prog_dly4 <= txcl_init_in_prog_dly3;
      end if;
    end if;
  end process;


-----------------------------------------------------------------------------
--  Start the TXD FSM
-----------------------------------------------------------------------------
  START_TX_DATA_FSM : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if set_start_txd_fsm = '1' then
        start_txd_fsm <= '1';
      else
        start_txd_fsm <= '0';
      end if;
    end if;
  end process;

-----------------------------------------------------------------------------
--  Delay the Enable for getting the End address
-----------------------------------------------------------------------------
  TXC_RD_END_ADDR_EN : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if set_txc_addr4_n = '1' then
        txc_rd_end    <= '1';
      else
        txc_rd_end    <= '0';
      end if;
      txc_rd_end_dly1 <= txc_rd_end;
    end if;
  end process;

-----------------------------------------------------------------------------
--  Store the end address
--    It will be used in Half Duplex mode to drop a packet if necessary
-----------------------------------------------------------------------------
  TXC_RD_END_ADDR : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        end_addr   <= (others => '0');
      else
        if txc_rd_end_dly1 = '1' then
          end_addr <= Tx_Client_TxC_2_Mem_Dout(c_TxD_addra_width -1 downto 0);
        else
          end_addr <= end_addr;
        end if;
      end if;
    end if;
  end process;


-----------------------------------------------------------------------------
--  Enable the memory
-----------------------------------------------------------------------------
  TXC_EN : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if set_txc_en = '1' then
        Tx_Client_TxC_2_Mem_En_int <= '1';
      else
        Tx_Client_TxC_2_Mem_En_int <= '0';
      end if;
    end if;
  end process;

  Tx_Client_TxC_2_Mem_En <= Tx_Client_TxC_2_Mem_En_int;

-----------------------------------------------------------------------------
--  Set the Write enable for memory writes
-----------------------------------------------------------------------------
  TXC_WR_EN : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if set_txc_wr = '1' then
        Tx_Client_TxC_2_Mem_We_int(0) <= '1';
      else
        Tx_Client_TxC_2_Mem_We_int(0) <= '0';
      end if;
    end if;
  end process;

  Tx_Client_TxC_2_Mem_We <= Tx_Client_TxC_2_Mem_We_int;

-----------------------------------------------------------------------------
--  Register the enable to align it with the Memory data
-----------------------------------------------------------------------------
  TXC_RD_EN : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      txc_wr_pntr_en <= set_txc_addr3;
    end if;
  end process;


  FIRST_RD_CMPLT : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        first_rd   <= '0';
      else
        if inc_txc_rd_addr = '1' then
          first_rd <= '1';
        else
          first_rd <= first_rd;
        end if;
      end if;
    end if;
  end process;

-----------------------------------------------------------------------------
--  TxC FIFO Data is captured on flop first to meet 2.5G timing requirement.
--  The FSM control signal is delated by 1 clock cycle to wait for the data to be available.
-----------------------------------------------------------------------------
  TXC_WRITE_POINTER_CAPTURE : process (tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txc_wr_pntr_2      <= (others => '0');
      else
        txc_wr_pntr_2      <= Tx_Client_TxC_2_Mem_Dout(c_TxC_addra_width -1 downto 0);
        if set_txc_addr3 = '1' and txc_wr_pntr_en = '1' then
          set_txc_addr3_d1 <= '1';
        else
          set_txc_addr3_d1 <= '0';
        end if;
      end if;
    end if;
  end process;

-----------------------------------------------------------------------------
--  TxC FIFO EMPTY Indicator
--    Compare the current TxC Rd Addr to the current TxC Wr Addr
-----------------------------------------------------------------------------
  TXC_WRITE_POINTER : process (tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txc_wr_pntr_1           <= (others => '0');
        txc_wr_pntr             <= (others => '0');
        compare_addr3_cmplt     <= '0';
      else
--------- if set_txc_addr3 = '1' and txc_wr_pntr_en = '1' then
        if set_txc_addr3_d1 = '1' then
          txc_wr_pntr_1         <= txc_wr_pntr_2;
          if txc_wr_pntr_1 = txc_wr_pntr_2 and compare_addr3_cmplt = '0' then
            txc_wr_pntr         <= txc_wr_pntr_1;
            compare_addr3_cmplt <= '1';
          else
            txc_wr_pntr         <= txc_wr_pntr;
            compare_addr3_cmplt <= '0';
          end if;
        else
          txc_wr_pntr_1         <= txc_wr_pntr_1;
          txc_wr_pntr           <= txc_wr_pntr;
          compare_addr3_cmplt   <= '0';
        end if;
      end if;
    end if;
  end process;

-----------------------------------------------------------------------------
--  Generate address that will get the End Address
-----------------------------------------------------------------------------
  TXC_RD_ADDR : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txc_mem_rd_addr       <= txc_min_rd_addr;
        txc_mem_rd_addr_0     <= txc_rd_addr5;
        txc_mem_rd_addr_1     <= txc_rd_addr6;
--  txc_rd_addr_cmp needs to lag one cnt because
--  it is incremented before the data is actually read
        txc_rd_addr_cmp       <= (others => '0');
      else
        if inc_txc_rd_addr = '1' and first_rd = '0' then
--  Initialize to start values
          txc_mem_rd_addr     <= txc_rd_addr5;
          txc_mem_rd_addr_0   <= txc_rd_addr6;
          txc_mem_rd_addr_1   <= txc_rd_addr7;
--  txc_rd_addr_cmp needs to lag one cnt because
--  it is incremented before the data is actually read
          txc_rd_addr_cmp     <= txc_min_rd_addr;
        elsif inc_txc_rd_addr = '1' and first_rd = '1' then
--  increment the address for the next packet
          if txc_mem_rd_addr = txc_max_rd_addr then
--  if the max address is reached, loop to address 0x4
            txc_mem_rd_addr   <= txc_mem_rd_addr_0;
            txc_mem_rd_addr_0 <= txc_mem_rd_addr_1;
            txc_mem_rd_addr_1 <= txc_rd_addr6;
            txc_rd_addr_cmp   <= txc_mem_rd_addr;
          else
--  otherwise just increment it
            txc_mem_rd_addr   <= txc_mem_rd_addr_0;
            txc_mem_rd_addr_0 <= txc_mem_rd_addr_1;
            txc_mem_rd_addr_1 <= std_logic_vector(unsigned(txc_mem_rd_addr_1) + 1);
            txc_rd_addr_cmp   <= txc_mem_rd_addr;
          end if;
        else                            -- Hold the current address until something changes
          txc_mem_rd_addr     <= txc_mem_rd_addr;
          txc_mem_rd_addr_0   <= txc_mem_rd_addr_0;
          txc_mem_rd_addr_1   <= txc_mem_rd_addr_1;
          txc_rd_addr_cmp     <= txc_rd_addr_cmp;
        end if;
      end if;
    end if;
  end process;


-----------------------------------------------------------------------------
--  Generate address mux fo memory
-----------------------------------------------------------------------------
  MEM_TXC_RD_ADDR : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if set_txc_addr4_n = '1' and first_rd = '0' and set_txc_wr = '0' then
-- Provide the address for the End of packet address
        Tx_Client_TxC_2_Mem_Addr_int <= txc_min_rd_addr;
      elsif set_txc_addr4_n = '1' and first_rd = '1' and set_txc_wr = '0' then
-- Provide the address for the End of packet address
        Tx_Client_TxC_2_Mem_Addr_int <= txc_mem_rd_addr;
      elsif set_txc_addr2 = '1' and set_txc_wr = '1' then
--Write the txc rd pointer
        Tx_Client_TxC_2_Mem_Addr_int <= txc_rd_addr2;
      elsif set_txc_addr3 = '1' and set_txc_wr = '0' then
--Read the txc wr pointer
        Tx_Client_TxC_2_Mem_Addr_int <= txc_rd_addr3;
      elsif set_txc_addr1 = '1' and set_txc_wr = '0' then
--  Read the TxD write pointer to monitor for an empty condition
        Tx_Client_TxC_2_Mem_Addr_int <= txc_rd_addr1;
      elsif set_txc_addr0 = '1' and set_txc_wr = '1' then
--  Write the current TxD Read Pointer while transmitting data
        Tx_Client_TxC_2_Mem_Addr_int <= txc_rd_addr0;
      else
        Tx_Client_TxC_2_Mem_Addr_int <= Tx_Client_TxC_2_Mem_Addr_int;
      end if;
    end if;
  end process;

  Tx_Client_TxC_2_Mem_Addr <= Tx_Client_TxC_2_Mem_Addr_int;

---------------------------------------------------------------------------
--  Write the TxC Rd Pointer to address 2 or
--    write the TxD Rd Pointer to address 0
--    Remove the lower 2 bits to align to a 32 bit word instead of a byte
---------------------------------------------------------------------------
  TXC_MEM_ADDR_PNTR : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if set_txc_addr2 = '1' then
--Address for data that is currently being transmitted
        Tx_Client_TxC_2_Mem_Din_int <= zeroes_txc & txc_rd_addr_cmp(c_TxC_addra_width -1 downto 0);
      elsif set_txc_addr0 = '1' then
        Tx_Client_TxC_2_Mem_Din_int <= zeroes_txd & txd_rd_addr(c_TxD_addra_width -1 downto 2);
      else
        Tx_Client_TxC_2_Mem_Din_int <= (others => '0');
      end if;
    end if;
  end process;

  Tx_Client_TxC_2_Mem_Din <= Tx_Client_TxC_2_Mem_Din_int;

-----------------------------------------------------------------------------
--  Transmit Client TX Control State Machine Combinatorial Logic
-----------------------------------------------------------------------------
    FSM_TXCLIENT_TXD_CMB : process (txd_rd_cs,tx_axis_mac_tready,
        start_txd_fsm,
        Tx_Client_TxD_2_Mem_Dout, txd_rd_addr,txc_rd_end,
        end_addr, phy_mode_enable, enabled_1588,
        tx_axis_mac_tready_dly, first_bytes)
    begin
        set_txd_vld      <= '0';
        clr_txd_vld      <= '0';
        set_txd_en       <= '0';
        inc_txd_rd_addr  <= '0';
        align_start_addr <= '0';
        set_txd_done     <= '0';
        mux_b3           <= '0';
        set_byte_en      <= '0';
        set_first_bytes  <= '0';
        txd_rd_ns        <= txd_rd_cs;

        case txd_rd_cs is
            when IDLE       =>
                if start_txd_fsm = '1' then
                    set_txd_en      <= '1';
                    if (enabled_1588 = '1') then
                        inc_txd_rd_addr <= '0';
                        set_first_bytes <= '0';
                        txd_rd_ns       <= GET_1588_CMD1;
                    else
                        inc_txd_rd_addr <= '1';
                        set_first_bytes <= '1';
                        txd_rd_ns       <= GET_B1;
                    end if;
                else
                    inc_txd_rd_addr <= '0';
                    set_txd_en      <= txc_rd_end;
                    txd_rd_ns       <= IDLE;
                end if;

            when GET_1588_CMD1 =>
                inc_txd_rd_addr   <= '1';
                set_txd_vld       <= '1'; 
                set_txd_en        <= '1';
                txd_rd_ns         <= GET_1588_CMD2;
            when GET_1588_CMD2 =>
                inc_txd_rd_addr   <= '1';
                set_txd_en        <= '1';
                txd_rd_ns         <= GET_1588_CMD3;
            when GET_1588_CMD3 =>
                inc_txd_rd_addr   <= '1';
                set_txd_en        <= '1';
                txd_rd_ns         <= GET_1588_CMD4;
            when GET_1588_CMD4 =>
                inc_txd_rd_addr   <= '1';
                set_txd_en        <= '1';
                txd_rd_ns         <= GET_1588_CMD5;
            when GET_1588_CMD5 =>
                inc_txd_rd_addr   <= '1';
                set_txd_en        <= '1';
                txd_rd_ns         <= GET_1588_CMD6;
            when GET_1588_CMD6 =>
                inc_txd_rd_addr   <= '1';
                set_txd_en        <= '1';
                txd_rd_ns         <= GET_1588_CMD7;
            when GET_1588_CMD7 =>
                inc_txd_rd_addr   <= '1';
                set_txd_en        <= '1';
                txd_rd_ns         <= GET_1588_CMD8;
            when GET_1588_CMD8 =>
                inc_txd_rd_addr   <= '1';
                set_txd_en        <= '1';
                set_first_bytes   <= '1';
                txd_rd_ns         <= GET_B1;

            when GET_B1     =>
                inc_txd_rd_addr   <= '1';
                set_txd_vld       <= '1'; --Start sending first data of payload
                set_txd_en        <= '1';
                txd_rd_ns         <= GET_B2;
            when GET_B2     =>
                inc_txd_rd_addr   <= '1';
                set_txd_en        <= '1';
                if (enabled_1588 = '0') then
                    set_byte_en       <= '1';
                end if;
                txd_rd_ns         <= GET_B3;
            when GET_B3     =>
                inc_txd_rd_addr   <= '1';
                set_txd_en        <= '1';
                txd_rd_ns         <= GET_B4;
                if (enabled_1588 = '1') then
                    set_byte_en       <= '1';
                end if;
            when GET_B4     =>
                txd_rd_ns         <= WAIT_TRDY2;
                if (enabled_1588 = '1') then
                    set_txd_en        <= '1';
                    inc_txd_rd_addr   <= '1';
                end if;
            when WAIT_TRDY2 =>
                if tx_axis_mac_tready = '1' and first_bytes = '0' and phy_mode_enable = '0' then
                    inc_txd_rd_addr <= '1'; --Continue reading payload data
                    set_txd_en      <= '1';
                    mux_b3          <= '1';
                    txd_rd_ns       <= WAIT_TRDY3;

                elsif tx_axis_mac_tready = '1' and first_bytes = '0' and phy_mode_enable = '1' then
                    inc_txd_rd_addr <= '0'; --Continue reading payload data
                    set_txd_en      <= '0';
                    mux_b3          <= '1';
                    txd_rd_ns       <= WAIT_TRDY3;

                else
                    inc_txd_rd_addr <= '0';
                    set_txd_en      <= '0';
                    mux_b3          <= '0';
                    txd_rd_ns       <= WAIT_TRDY2;
                end if;

            when WAIT_TRDY3 =>
                if tx_axis_mac_tready = '1' then
                    inc_txd_rd_addr <= '1'; --Continue reading payload data
                    set_txd_en      <= '1';
                    txd_rd_ns       <= CHECK_DONE;
                else
                    inc_txd_rd_addr <= '0';
                    set_txd_en      <= '0';
                    txd_rd_ns       <= WAIT_TRDY3;
                end if;

            when CHECK_DONE =>
                if tx_axis_mac_tready = '1' then
--  The end addreess read from the memory is always one byte before
--  the actual end of the packet to allow tlast to be asserted correctly

--  On the write side of the BRAM, the end_addr has been set such that the
--  at strobes at TLAST reflect the last byte of data minus 1
--    case axi_str_txd_tstrb_dly0 is
--      when "1111" => end_addr_byte_offset <= "11";
--      when "0111" => end_addr_byte_offset <= "10";
--      when "0011" => end_addr_byte_offset <= "01";
--      when others => end_addr_byte_offset <= "00";
--    end case;
--
--  The BRAM parity bits are not used with AXI-S CORE Gen
--
                    if end_addr = txd_rd_addr then
--Last byte of payload data is one byte after end_address
                        if txd_rd_addr(1) = '1' and txd_rd_addr (0) = '1' then
--  By incrementing the address one, it will be 32 bit aligned
--  which is the starting address of the next packet
                            align_start_addr <= '0';
                            inc_txd_rd_addr  <= '1';
                        else
--  Align address to 32 bits because it ended non aligned
--    The next 32 bit aligned address will be the start
--    of the next payload data
--  Do not increment the address since it is getting aligned
                            align_start_addr <= '1';
                            inc_txd_rd_addr  <= '0';
                        end if;
                        if phy_mode_enable = '0' then
                            clr_txd_vld      <= '0';
                            set_txd_en       <= '0';
                            set_txd_done     <= '0';
                            txd_rd_ns        <= WAIT_LAST;
                        elsif phy_mode_enable = '1' then
                            clr_txd_vld      <= '1';
                            set_txd_en       <= '0';
                            set_txd_done     <= '1';
                            txd_rd_ns        <= IDLE;
                        end if;
                    else
                        inc_txd_rd_addr    <= '1'; --set addr to get next data
                        set_txd_en         <= '1';
                        set_txd_done       <= '0';
                        align_start_addr   <= '0';
                        txd_rd_ns          <= CHECK_DONE;
                    end if;
                else
                    inc_txd_rd_addr      <= '0';
                    set_txd_en           <= '0';
                    set_txd_done         <= '0';
                    align_start_addr     <= '0';
                    txd_rd_ns            <= CHECK_DONE;
                end if;

            when WAIT_LAST =>
--  Need to wait one tready clock cycle before transitioning to IDLE
--    This will allow the last Tx Byte through and set TLAST accordingly
                clr_txd_vld     <= '1';
                inc_txd_rd_addr <= '0';
                set_txd_en      <= '0';
                set_txd_done    <= '1';
                txd_rd_ns       <= IDLE;

            when others =>
                txd_rd_ns <= IDLE;

        end case;
    end process;

-----------------------------------------------------------------------------
--  Transmit Client TX Control State Machine Sequencer
-----------------------------------------------------------------------------
    FSM_TXCLIENT_TXD_SEQ : process (tx_axi_clk)
    begin
        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd_rd_cs <= IDLE;
                set_txd_vld_1       <= '0';
                set_txd_vld_2       <= '0';
            else
                txd_rd_cs <= txd_rd_ns;
                set_txd_vld_1       <= set_txd_vld and enabled_1588;
                set_txd_vld_2       <= set_txd_vld_1 and enabled_1588;
            end if;
        end if;
    end process;


-----------------------------------------------------------------------------
--  Transmit Client TX Complete Signal
-----------------------------------------------------------------------------
    TX_COMPLETE_INDICATOR : process (tx_axi_clk)
    begin
        if rising_edge(tx_axi_clk) then
            if set_txd_done = '1' then
                tx_cmplt <= '1';
            else
                tx_cmplt <= '0';
            end if;
        end if;
    end process;

-----------------------------------------------------------------------------
--  Set byte enable pipeline to use individual bits to store the BRAM data
--  as it is read.  Then use the stored data to send to the MAC when
--  appropriate.
-----------------------------------------------------------------------------
    BX_EN_PIPE : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if set_byte_en = '1' then
                set_byte_en_pipe(0) <= '1';
            else
                set_byte_en_pipe(0) <= '0';
            end if;
            set_byte_en_pipe(1)   <= set_byte_en_pipe(0);
        end if;
    end process;


-----------------------------------------------------------------------------
--  Store Byte 1 data so it can be muxed to txd on each packets first
--  tx_axis_mac_tready assertion
-----------------------------------------------------------------------------
    TXD_BYTE1 : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd_1   <= (others => '0');
            else
                if set_byte_en = '1' then
                    txd_1 <= Tx_Client_TxD_2_Mem_Dout(C_CLIENT_WIDTH-1 downto 0);
                else
                    txd_1 <= txd_1;
                end if;
            end if;
        end if;
    end process;


-----------------------------------------------------------------------------
--  Store Byte 2 data so it can be muxed to txd on each packets second
--  tx_axis_mac_tready assertion
-----------------------------------------------------------------------------
    TXD_BYTE2 : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd_2   <= (others => '0');
            else
                if set_byte_en_pipe(0) = '1' then
                    txd_2 <= Tx_Client_TxD_2_Mem_Dout(C_CLIENT_WIDTH-1 downto 0);
                else
                    txd_2 <= txd_2;
                end if;

            end if;
        end if;
    end process;


-----------------------------------------------------------------------------
--  Store Byte 3 data so it can be muxed to txd on each packets third
--  tx_axis_mac_tready assertion
-----------------------------------------------------------------------------
    TXD_BYTE3 : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd_3   <= (others => '0');
            else
                if set_byte_en_pipe(1) = '1' then
                    txd_3 <= Tx_Client_TxD_2_Mem_Dout(C_CLIENT_WIDTH-1 downto 0);
                else
                    txd_3 <= txd_3;
                end if;

            end if;
        end if;
    end process;


-----------------------------------------------------------------------------
--  Use this delay to mux in the stored first bytes of data for each packet
-----------------------------------------------------------------------------
    TX_ACK_DELAY : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then

            if tx_axis_mac_tready = '1' then
                tx_axis_mac_tready_dly <= '1';
            else
                tx_axis_mac_tready_dly <= '0';
            end if;
        end if;

    end process;

-----------------------------------------------------------------------------
--  TxD Read Memory Enable - only enable memory when needed
-----------------------------------------------------------------------------
    TXD_MEM_EN : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if set_txd_en = '1' then
                Tx_Client_TxD_2_Mem_En_int <= '1';
            else
                Tx_Client_TxD_2_Mem_En_int <= '0';
            end if;
        end if;
    end process;

    Tx_Client_TxD_2_Mem_En <= Tx_Client_TxD_2_Mem_En_int;

-----------------------------------------------------------------------------
--  TxD Memory Write Enable bit is never written to
-----------------------------------------------------------------------------
    Tx_Client_TxD_2_Mem_We(0) <= '0';

-----------------------------------------------------------------------------
--  Get Lower 2 bits for case statement below
-----------------------------------------------------------------------------
    txd_rd_addr_1_0 <= txd_rd_addr(1 downto 0); -- for case statement below

-----------------------------------------------------------------------------
--  Set the address to be 32 bit aligned for readjustment at the end of
--    the packet
-----------------------------------------------------------------------------
  txd_rd_addr_aligned <= txd_rd_addr(c_TxD_addra_width -1 downto 2) & "00";

-----------------------------------------------------------------------------
--  Generate the TxD Memory Read Address
-----------------------------------------------------------------------------
      TXD_MEM_RD_ADDR : process(tx_axi_clk)
      begin
  
        if rising_edge(tx_axi_clk) then
          if reset2tx_client = '1' then
            txd_rd_addr     <= (others => '0');
          else
--  the end of the packet was reached, so adjust the Rd Addr
--    to be 32bit aligned if needed
            if align_start_addr = '1' then
              case txd_rd_addr_1_0 is
                when "00" | "01" | "10" => --  | "11" =>
-- packet ended on a non 32bit aligned address, so adjust it
                  txd_rd_addr <= std_logic_vector(unsigned(txd_rd_addr_aligned) + 4);
                when  others =>
-- packet ended on a 32bit aligned address, so do not change
                  txd_rd_addr <= txd_rd_addr;
              end case;
            else
--  increment to next address
              if inc_txd_rd_addr = '1' then
                txd_rd_addr <= std_logic_vector(unsigned(txd_rd_addr) + 1);
              else
                txd_rd_addr <= txd_rd_addr;
              end if;
            end if;
          end if;
        end if;
      end process;

        Tx_Client_TxD_2_Mem_Addr <= txd_rd_addr;


---------------------------------------------------------------------------
--  Force and update the BRAM with the rd_pntr_addr every ~512 bytes
---------------------------------------------------------------------------
    BRAM_UPDATE : process(tx_axi_clk)
    begin
        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' or set_txd_done = '1' then
                update_bram_cnt   <= (others => '0');
            else
                if update_bram_cnt(9) = '1' and inc_txd_rd_addr = '1' then
                    update_bram_cnt <= ('0' & update_bram_cnt(8 downto 0)) + 1;
                elsif inc_txd_rd_addr = '1' then
                    update_bram_cnt <= update_bram_cnt + 1;
                else
                    update_bram_cnt <= update_bram_cnt;
                end if;
            end if;
        end if;
    end process;


---------------------------------------------------------------------------
--  Use this signal to dis-allow a transition to the WAIT_TRDY3 state of
--  the FSM_TXCLIENT_TXD_CMB FSM when in the WAIT_TRDY2 state
---------------------------------------------------------------------------
        SET_FIRST_BYTE_FILTER : process (tx_axi_clk)
        begin
          if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' or (tx_axis_mac_tready = '0' and tx_axis_mac_tready_dly = '1') then
              first_bytes   <= '0';
            else
              if set_first_bytes = '1' then
                first_bytes <= '1';
              else
                first_bytes <= first_bytes;
              end if;
            end if;
          end if;
        end process;


-----------------------------------------------------------------------------
--  Mux the Memory data to the Tx Client Interface when appropriate
--    1. Mux the first byte
--    2. Mux the second byte at the rising edge of the first tready of the packet
--    3. Mux the third byte at the second tready of the packet
--    4. Mux the fourth byte at the third tready of the packet
--    5. Mux the remaining bytes
-----------------------------------------------------------------------------
    TXD_MEM_DATA : process (tx_axi_clk)
    begin
        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd   <= (others => '0');
            else
                if set_txd_vld = '1' or set_txd_vld_1 = '1'  or set_txd_vld_2 = '1'then
                    txd <= Tx_Client_TxD_2_Mem_Dout(C_CLIENT_WIDTH-1 downto 0); --load first byte and hold until ack
                elsif tx_axis_mac_tready = '1' and tx_axis_mac_tready_dly = '0' and first_bytes = '1' then
                    txd <= txd_1;
                elsif tx_axis_mac_tready = '0' and tx_axis_mac_tready_dly = '1' and first_bytes = '1' then
                    txd <= txd_2;
                elsif tx_axis_mac_tready = '1' and tx_axis_mac_tready_dly = '1' and first_bytes = '1' then
                    txd <= txd_2;
                elsif mux_b3 = '1' then
                    txd <= txd_3;
                elsif tx_axis_mac_tready = '1' then
                    txd <= Tx_Client_TxD_2_Mem_Dout(C_CLIENT_WIDTH -1 downto 0); --remaining bytes
                else
                    txd <= txd;
                end if;
            end if;
        end if;
    end process;

    tx_axis_mac_tdata <= txd;

-----------------------------------------------------------------------------
--  Assert Transmit Data Valid for the duration of a transmitted packet
-----------------------------------------------------------------------------
    SET_TX_DATA_VALID : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd_vld   <= '0';
            else
                if tx_axis_mac_tready = '1' and tx_axis_mac_tlast_int = '1' then
                    txd_vld <= '0';
                elsif set_txd_vld = '1' then
                    txd_vld <= '1';
                else
                    txd_vld <= txd_vld;
                end if;
            end if;
        end if;
    end process;

    tx_axis_mac_tvalid <= txd_vld;

-----------------------------------------------------------------------------
--  Assert Transmit Data LAST to end the packet
-----------------------------------------------------------------------------
    SET_TLAST : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                tx_axis_mac_tlast_int   <= '0';
            elsif tx_axis_mac_tready = '1' then
                if clr_txd_vld = '1' then
                    tx_axis_mac_tlast_int <= '1';
                else
                    tx_axis_mac_tlast_int <= '0';
                end if;
            else
                tx_axis_mac_tlast_int   <= tx_axis_mac_tlast_int;
            end if;
        end if;
    end process;

    tx_axis_mac_tlast <= tx_axis_mac_tlast_int;

-----------------------------------------------------------------------------
--  Register the Enable to align it with the TxC Memory Dout Write pointer
--    Hold the enable from the start of the packet to the end of the packet
-----------------------------------------------------------------------------
    TXD_WR_POINTER_EN : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' or (txd_wr_pntr_en = '1' and tx_axis_mac_tready = '1') then
                txd_wr_pntr_en <= '0';
            elsif set_txc_addr0 = '1' then
                txd_wr_pntr_en <= '1';
            else
                txd_wr_pntr_en <= txd_wr_pntr_en;
            end if;
        end if;
    end process;

end rtl;


-------------------------------------------------------------------------------
-- tx_emac_if_2g5 - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename: tx_emac_if_2g5.vhd
-- Version: v1.00a
-- Description: top level of embedded ip Ethernet MAC interface
--
-- VHDL-Standard: VHDL'93
-------------------------------------------------------------------------------
-- Structure: This section shows the hierarchical structure of axi_ethernet.
--
-- axi_ethernet.vhd
-- axi_ethernt_soft_temac_wrap.vhd
-- axi_lite_ipif.vhd
-- embedded_top.vhd
-- tx_if.vhd
-- tx_axistream_if.vhd
-- tx_mem_if
-- -> tx_emac_if_2g5.vhd
--
-------------------------------------------------------------------------------
-- Author: vineelc
--
-- vineelc 11/27/23
-- ^^^^^^
-- - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
-- active low signals: "*_n"
-- clock signals: "clk", "clk_div#", "clk_#x"
-- reset signals: "rst", "rst_n"
-- generics: "C_*"
-- user defined types: "*_TYPE"
-- state machine next state: "*_ns"
-- state machine current state: "*_cs"
-- combinatorial signals: "*_com"
-- pipelined or register delay signals: "*_d#"
-- counter signals: "*cnt*"
-- clock enable signals: "*_ce"
-- internal version of output port "*_i"
-- device pins: "*_pin"
-- ports: - Names begin with Uppercase
-- processes: "*_PROCESS"
-- component instantiations: "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tx_if_pack.all;


-------------------------------------------------------------------------------
-- Entity Section
-------------------------------------------------------------------------------

entity tx_emac_if_2g5 is
  generic (
    C_FAMILY            : string                   := "virtex6";
    C_HALFDUP           : integer range 0 to 1     := 0;
    C_TXMEM             : integer                  := 4096;
    C_TXCSUM            : integer range 0 to 2     := 0;
    C_ENABLE_1588       : integer                  := 0;

-- Read Port - AXI Stream TxData
    c_TxD_write_width_a : integer range 0 to 18    := 9;
    c_TxD_read_width_a  : integer range 0 to 18    := 9;
    c_TxD_write_depth_a : integer range 0 to 32768 := 4096;
    c_TxD_read_depth_a  : integer range 0 to 32768 := 4096;
    c_TxD_addra_width   : integer range 0 to 15    := 10;
    c_TxD_wea_width     : integer range 0 to 2     := 2;

-- Read Port - AXI Stream TxControl
    c_TxC_write_width_a : integer range 36 to 36   := 36;
    c_TxC_read_width_a  : integer range 36 to 36   := 36;
    c_TxC_write_depth_a : integer range 0 to 1024  := 1024;
    c_TxC_read_depth_a  : integer range 0 to 1024  := 1024;
    c_TxC_addra_width   : integer range 0 to 10    := 10;
    c_TxC_wea_width     : integer range 0 to 1     := 1;

    c_TxD_addrb_width   : integer range 0 to 13    := 10;

    C_CLIENT_WIDTH      : integer                  := 8
    );
  port (
--Transmit Memory Read Interface
-- ** WARNING ** WARNING ** WARNING **
--  For MII,GMII, RGMI, 1000Base-X and pcs/pma SGMII this is an accurate indicator
--  However for V6 Hard SGMII it is always tied to '0' for all speeds
    tx_client_10_100         : in  std_logic; --  Tx Client CE Toggles Indicator

-- Read Port - AXI Stream TxData
    reset2tx_client          : in  std_logic; --  reset
    Tx_Client_TxD_2_Mem_Din  : out std_logic_vector (c_TxD_write_width_a-1 downto 0); --  Tx AXI-Stream Data to Memory Wr Din
    Tx_Client_TxD_2_Mem_Addr : out std_logic_vector (c_TxD_addra_width-1 downto 0  ); --  Tx AXI-Stream Data to Memory Wr Addr
    Tx_Client_TxD_2_Mem_En   : out std_logic; --  Tx AXI-Stream Data to Memory Enable
    Tx_Client_TxD_2_Mem_We   : out std_logic_vector (c_TxD_wea_width-1 downto 0    ); --  Tx AXI-Stream Data to Memory Wr En
    Tx_Client_TxD_2_Mem_Dout : in  std_logic_vector (c_TxD_read_width_a-1 downto 0 ); --  Tx AXI-Stream Data to Memory Not Used

-- Read Port - AXI Stream TxControl
    reset2axi_str_txd        : in  std_logic; --  reset
    Tx_Client_TxC_2_Mem_Din  : out std_logic_vector (c_TxC_write_width_a-1 downto 0); --  Tx AXI-Stream Control to Memory Wr Din
    Tx_Client_TxC_2_Mem_Addr : out std_logic_vector (c_TxC_addra_width-1 downto 0  ); --  Tx AXI-Stream Control to Memory Wr Addr
    Tx_Client_TxC_2_Mem_En   : out std_logic; --  Tx AXI-Stream Control to Memory Enable
    Tx_Client_TxC_2_Mem_We   : out std_logic_vector (c_TxC_wea_width-1 downto 0    ); --  Tx AXI-Stream Control to Memory Wr En
    Tx_Client_TxC_2_Mem_Dout : in  std_logic_vector (c_TxC_read_width_a-1 downto 0 ); --  Tx AXI-Stream Control to Memory Full Flag

--  Tx AXI-S Interface
    tx_axi_clk               : in  std_logic; --  Tx AXI-Stream clock in
    tx_reset_out             : in  std_logic; --  take to reset combiner
    tx_axis_mac_tdata        : out std_logic_vector (C_CLIENT_WIDTH - 1 downto 0   ); --  Tx AXI-Stream data
    tx_axis_mac_tvalid       : out std_logic; --  Tx AXI-Stream valid
    tx_axis_mac_tlast        : out std_logic; --  Tx AXI-Stream last
    tx_axis_mac_tuser        : out std_logic; -- this is always driven low since an underflow cannot occur
    tx_axis_mac_tready       : in  std_logic; --  Tx AXI-Stream ready in from TEMAC
    tx_collision             : in  std_logic; --  collision not used
    tx_retransmit            : in  std_logic; -- retransmit not used


    tx_cmplt                 : out std_logic; -- transmit is complete indicator

    tx_init_in_prog_cross    : in  std_logic        --  Tx is Initializing after a reset
    );

end tx_emac_if_2g5;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of tx_emac_if_2g5 is

    type TXC_RD_FSM_TYPE is (
    GET_TXC_WR_PNTR,
    GET_END_PNTR,
    SET_TXCRD_PNTR,
    GET_TXDWR_PNTR,
    SET_TXDRD_PNTR,
    WAIT_TXD_DONE,
    GET_ADDR3,
    WAIT_ADDR3_PNTR);

    signal txc_rd_cs, txc_rd_ns : TXC_RD_FSM_TYPE;

    type TXD_RD_FSM_TYPE is (
    IDLE,
    GET_B1,
    WAIT_TRDY,
    STREAM_DATA,
    WAIT_LAST);

    signal txd_rd_cs, txd_rd_ns : TXD_RD_FSM_TYPE;

    signal enable_1588_val     : std_logic_vector(2 downto 0) := (others => '0'); 
    signal enabled_1588        : std_logic;
    signal set_txc_addr0       : std_logic;
    signal set_txc_addr1       : std_logic;
    signal set_txc_addr2       : std_logic;
    signal set_txc_addr3       : std_logic;
    signal set_txc_addr3_d1    : std_logic;
    signal txc_addr3_en        : std_logic;
    signal set_txc_addr4_n     : std_logic;
    signal set_txc_wr          : std_logic;
    signal set_txc_en          : std_logic;
    signal txc_wr_pntr_en      : std_logic;
    signal set_start_txd_fsm   : std_logic;
    signal start_txd_fsm       : std_logic;
    signal inc_txc_rd_addr     : std_logic;
    signal first_rd            : std_logic;
    signal txc_wr_pntr_1       : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_wr_pntr_2       : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_wr_pntr         : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal compare_addr3_cmplt : std_logic;

    signal Tx_Client_TxC_2_Mem_Addr_int : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_mem_rd_addr              : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr_cmp              : std_logic_vector(c_TxC_addra_width -1 downto 0);

    signal end_addr                    : std_logic_vector(c_TxD_addra_width -1 downto 0);
    signal txc_rd_end                  : std_logic;
    signal txc_rd_end_dly1             : std_logic;
    signal Tx_Client_TxC_2_Mem_En_int  : std_logic;
    signal Tx_Client_TxC_2_Mem_We_int  : std_logic_vector(c_TxC_wea_width-1 downto 0);
    signal Tx_Client_TxC_2_Mem_Din_int : std_logic_vector(c_TxC_write_width_a -1 downto 0);

    signal set_txd_vld            : std_logic;
    signal clr_txd_vld            : std_logic;
	signal clr_txd_vld_d1         : std_logic;
    signal set_txd_en             : std_logic;
    signal inc_txd_rd_addr        : std_logic;
    signal txd_rd_addr            : std_logic_vector(c_TxD_addra_width -1 downto 0);
    signal txd_rd_addr_1_0        : std_logic_vector(1 downto 0);
    signal txd_rd_addr_aligned    : std_logic_vector(c_TxD_addra_width -1 downto 0);

    signal align_start_addr           : std_logic;
    signal set_txd_done               : std_logic;
    signal Tx_Client_TxD_2_Mem_En_int : std_logic;
    signal txd                        : std_logic_vector(C_CLIENT_WIDTH-1 downto 0);
    signal txd_vld                    : std_logic;

    signal txc_min_rd_addr : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_max_rd_addr : std_logic_vector(c_TxC_addra_width -1 downto 0);

    signal txc_rd_addr0 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr1 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr2 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr3 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr5 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr6 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_rd_addr7 : std_logic_vector(c_TxC_addra_width -1 downto 0);

    signal txc_mem_rd_addr_0 : std_logic_vector(c_TxC_addra_width -1 downto 0);
    signal txc_mem_rd_addr_1 : std_logic_vector(c_TxC_addra_width -1 downto 0);

    signal txd_pipe : std_logic_vector(C_CLIENT_WIDTH-1 downto 0);


    constant zeroes_txc : std_logic_vector(c_TxC_read_width_a -1 downto c_TxC_addra_width)    := (others => '0');
    constant zeroes_txd : std_logic_vector(c_TxC_read_width_a -1 downto c_TxD_addra_width -2) := (others => '0');

    signal txcl_init_in_prog_dly1 : std_logic;
    signal txcl_init_in_prog_dly2 : std_logic;
    signal txcl_init_in_prog_dly3 : std_logic;
    signal txcl_init_in_prog_dly4 : std_logic;

    signal update_bram_cnt : unsigned(9 downto 0);

    signal tx_axis_mac_tready_dly : std_logic;

    signal tx_axis_mac_tlast_int : std_logic;

    signal load_tx_pipe          : std_logic;
	signal flush_tx_pipe         : std_logic;


    signal phy_mode_enable : std_logic;

begin

    tx_axis_mac_tuser <= '0';

    Tx_Client_TxD_2_Mem_Din <= (others => '0');

    phy_mode_enable <= tx_client_10_100;

    enable_1588_val <= std_logic_vector(to_unsigned(C_ENABLE_1588, enable_1588_val'length));
    enabled_1588 <= '1' when ((enable_1588_val(1) = '1' and enable_1588_val(0) = '0') or (enable_1588_val(1) = '0' and enable_1588_val(0) = '1')) 
                    else '0';

-----------------------------------------------------------------------------
--  Create the full and empty comparison values for the S6 and V6 since
--  1 S6 BRAM = 1/2 V6 BRAM
-----------------------------------------------------------------------------
    GEN_TXC_MIN_MAX_RD_FLAG : for i in (c_TxC_addra_width - 1) downto 0 generate
        txc_min_rd_addr(i) <= '1' when (i = 2)                   else '0';
        txc_max_rd_addr(i) <= '0' when (i = 0 or i = 1)          else '1';
        txc_rd_addr0(i)    <= '0';
        txc_rd_addr1(i)    <= '1' when (i = 0)                   else '0';
        txc_rd_addr2(i)    <= '1' when (i = 1)                   else '0';
        txc_rd_addr3(i)    <= '1' when (i = 0 or i = 1)          else '0';
        txc_rd_addr5(i)    <= '1' when (i = 0 or i = 2)          else '0';
        txc_rd_addr6(i)    <= '1' when (i = 1 or i = 2)          else '0';
        txc_rd_addr7(i)    <= '1' when (i = 0 or i = 1 or i = 2) else '0';

    end generate GEN_TXC_MIN_MAX_RD_FLAG;

-----------------------------------------------------------------------------
--  Transmit Client TX Control State Machine Combinatorial Logic
-----------------------------------------------------------------------------
    FSM_TXCLIENT_TXC_CMB : process (txc_rd_cs,tx_axis_mac_tready,
      clr_txd_vld,txc_rd_addr_cmp,
      txcl_init_in_prog_dly4,compare_addr3_cmplt,txc_wr_pntr,
      update_bram_cnt)
    begin
        set_txc_addr0     <= '0';
        set_txc_addr1     <= '0';
        set_txc_addr2     <= '0';
        set_txc_addr3     <= '0';
        set_txc_addr4_n   <= '0';
        set_txc_wr        <= '0';
        set_txc_en        <= '0';
        set_start_txd_fsm <= '0';
        inc_txc_rd_addr   <= '0';

        case txc_rd_cs is
            when GET_TXC_WR_PNTR =>
                if txcl_init_in_prog_dly4 = '0' and compare_addr3_cmplt = '1' and txc_rd_addr_cmp /= txc_wr_pntr then
                    set_txc_addr3     <= '0';
                    set_txc_addr4_n   <= '1'; -- Read TxC Addr 0x4 - 0xn
                    set_txc_en        <= '1';
                    inc_txc_rd_addr   <= '1';
                    txc_rd_ns         <= GET_END_PNTR;
                else
                    set_txc_addr3     <= '1'; -- Read TxC Addr 0x3 (TxC Empty)
                    set_txc_addr4_n   <= '0';
                    set_txc_en        <= '1';
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= GET_TXC_WR_PNTR;
                end if;
            when GET_END_PNTR    =>
                set_txc_addr2       <= '1'; -- Write TxC Addr 0x2
                set_txc_wr          <= '1';
                set_txc_en          <= '1';
                txc_rd_ns           <= SET_TXCRD_PNTR;
            when SET_TXCRD_PNTR  =>
                set_txc_addr1       <= '1'; -- Read TxC Addr 0x1
                set_txc_en          <= '1';
                txc_rd_ns           <= GET_TXDWR_PNTR;
            when GET_TXDWR_PNTR  =>
                set_txc_addr0       <= '1'; -- Write TxC Addr 0x0
                set_txc_wr          <= '1';
                set_txc_en          <= '1';
                txc_rd_ns           <= SET_TXDRD_PNTR;
            when SET_TXDRD_PNTR  =>
                set_txc_addr0       <= '0';
                set_txc_wr          <= '0';
                set_txc_en          <= '0';
                set_start_txd_fsm   <= '1';
                txc_rd_ns           <= WAIT_TXD_DONE;
            when WAIT_TXD_DONE   =>
                if tx_axis_mac_tready = '1' and clr_txd_vld = '0' then
                    if update_bram_cnt(9) = '1' then  --Update the TxC BRAM with the current rd_addr_addr
                        set_txc_addr0   <= '1'; -- Write TxC Addr 0x0
                        set_txc_addr3   <= '0';
                        set_txc_wr      <= '1';
                        set_txc_en      <= '1';
                        inc_txc_rd_addr <= '0';
                        txc_rd_ns       <= WAIT_TXD_DONE;
                    else
                        set_txc_addr0   <= '0'; -- Write TxC Addr 0x0
                        set_txc_addr3   <= '0';
                        set_txc_wr      <= '0';
                        set_txc_en      <= '0';
                        inc_txc_rd_addr <= '0';
                        txc_rd_ns       <= WAIT_TXD_DONE;
                    end if;
                elsif tx_axis_mac_tready = '1' and clr_txd_vld = '1' then
                    set_txc_addr0     <= '1';
                    set_txc_addr3     <= '0';
                    set_txc_wr        <= '1';
                    set_txc_en        <= '1'; --write the last rd_rntr_addr for this packet
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= GET_ADDR3;
                else
                    set_txc_addr0     <= '0';
                    set_txc_addr3     <= '0'; --do nothing
                    set_txc_wr        <= '0';
                    set_txc_en        <= '0';
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= WAIT_TXD_DONE;
                end if;
            when GET_ADDR3       =>
                if tx_axis_mac_tready = '1' then
                    set_txc_addr0     <= '0';
                    set_txc_addr3     <= '1';
                    set_txc_wr        <= '0';
                    set_txc_en        <= '1'; --get ready for the next packet - addr0x4-0xn
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= WAIT_ADDR3_PNTR;
                else
                    set_txc_addr0     <= '0';
                    set_txc_addr3     <= '0';
                    set_txc_wr        <= '0';
                    set_txc_en        <= '0';
                    inc_txc_rd_addr   <= '0';
                    txc_rd_ns         <= GET_ADDR3;
                end if;
            when WAIT_ADDR3_PNTR =>
                set_txc_addr0       <= '0';
                set_txc_addr3       <= '1';
                set_txc_wr          <= '0';
                set_txc_en          <= '1';
                inc_txc_rd_addr     <= '0';
                txc_rd_ns           <= GET_TXC_WR_PNTR;
            when others          =>
                txc_rd_ns           <= GET_TXC_WR_PNTR;
        end case;
    end process;

-----------------------------------------------------------------------------
--  Transmit Client TX Control State Machine Sequencer
-----------------------------------------------------------------------------
  FSM_TXCLIENT_TXC_SEQ : process (tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txc_rd_cs <= GET_TXC_WR_PNTR;
      else
        txc_rd_cs <= txc_rd_ns;
      end if;
    end if;
  end process;

---------------------------------------------------------------------------
--  Delay the indicator to ensure the memory has had enough time to update
---------------------------------------------------------------------------
  TXCL_INIT_INDICATOR_DLY : process (tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txcl_init_in_prog_dly1 <= '1';
        txcl_init_in_prog_dly2 <= '1';
        txcl_init_in_prog_dly3 <= '1';
        txcl_init_in_prog_dly4 <= '1';
      else
        txcl_init_in_prog_dly1 <= tx_init_in_prog_cross;
        txcl_init_in_prog_dly2 <= txcl_init_in_prog_dly1;
        txcl_init_in_prog_dly3 <= txcl_init_in_prog_dly2;
        txcl_init_in_prog_dly4 <= txcl_init_in_prog_dly3;
      end if;
    end if;
  end process;


-----------------------------------------------------------------------------
--  Start the TXD FSM
-----------------------------------------------------------------------------
  START_TX_DATA_FSM : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if set_start_txd_fsm = '1' then
        start_txd_fsm <= '1';
      else
        start_txd_fsm <= '0';
      end if;
    end if;
  end process;

-----------------------------------------------------------------------------
--  Delay the Enable for getting the End address
-----------------------------------------------------------------------------
  TXC_RD_END_ADDR_EN : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if set_txc_addr4_n = '1' then
        txc_rd_end    <= '1';
      else
        txc_rd_end    <= '0';
      end if;
      txc_rd_end_dly1 <= txc_rd_end;
    end if;
  end process;

-----------------------------------------------------------------------------
--  Store the end address
--    It will be used in Half Duplex mode to drop a packet if necessary
-----------------------------------------------------------------------------
  TXC_RD_END_ADDR : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        end_addr   <= (others => '0');
      else
        if txc_rd_end_dly1 = '1' then
          end_addr <= Tx_Client_TxC_2_Mem_Dout(c_TxD_addra_width -1 downto 0);
        else
          end_addr <= end_addr;
        end if;
      end if;
    end if;
  end process;


-----------------------------------------------------------------------------
--  Enable the memory
-----------------------------------------------------------------------------
  TXC_EN : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if set_txc_en = '1' then
        Tx_Client_TxC_2_Mem_En_int <= '1';
      else
        Tx_Client_TxC_2_Mem_En_int <= '0';
      end if;
    end if;
  end process;

  Tx_Client_TxC_2_Mem_En <= Tx_Client_TxC_2_Mem_En_int;

-----------------------------------------------------------------------------
--  Set the Write enable for memory writes
-----------------------------------------------------------------------------
  TXC_WR_EN : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if set_txc_wr = '1' then
        Tx_Client_TxC_2_Mem_We_int(0) <= '1';
      else
        Tx_Client_TxC_2_Mem_We_int(0) <= '0';
      end if;
    end if;
  end process;

  Tx_Client_TxC_2_Mem_We <= Tx_Client_TxC_2_Mem_We_int;

-----------------------------------------------------------------------------
--  Register the enable to align it with the Memory data
-----------------------------------------------------------------------------
  TXC_RD_EN : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      txc_wr_pntr_en <= set_txc_addr3;
    end if;
  end process;


  FIRST_RD_CMPLT : process(tx_axi_clk)
  begin

    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        first_rd   <= '0';
      else
        if inc_txc_rd_addr = '1' then
          first_rd <= '1';
        else
          first_rd <= first_rd;
        end if;
      end if;
    end if;
  end process;

-----------------------------------------------------------------------------
--  TxC FIFO Data is captured on flop first to meet 2.5G timing requirement.
--  The FSM control signal is delated by 1 clock cycle to wait for the data to be available.
-----------------------------------------------------------------------------
  TXC_WRITE_POINTER_CAPTURE : process (tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txc_wr_pntr_2      <= (others => '0');
      else
        txc_wr_pntr_2      <= Tx_Client_TxC_2_Mem_Dout(c_TxC_addra_width -1 downto 0);
        if set_txc_addr3 = '1' and txc_wr_pntr_en = '1' then
          set_txc_addr3_d1 <= '1';
        else
          set_txc_addr3_d1 <= '0';
        end if;
      end if;
    end if;
  end process;

-----------------------------------------------------------------------------
--  TxC FIFO EMPTY Indicator
--    Compare the current TxC Rd Addr to the current TxC Wr Addr
-----------------------------------------------------------------------------
  TXC_WRITE_POINTER : process (tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txc_wr_pntr_1           <= (others => '0');
        txc_wr_pntr             <= (others => '0');
        compare_addr3_cmplt     <= '0';
      else
--------- if set_txc_addr3 = '1' and txc_wr_pntr_en = '1' then
        if set_txc_addr3_d1 = '1' then
          txc_wr_pntr_1         <= txc_wr_pntr_2;
          if txc_wr_pntr_1 = txc_wr_pntr_2 and compare_addr3_cmplt = '0' then
            txc_wr_pntr         <= txc_wr_pntr_1;
            compare_addr3_cmplt <= '1';
          else
            txc_wr_pntr         <= txc_wr_pntr;
            compare_addr3_cmplt <= '0';
          end if;
        else
          txc_wr_pntr_1         <= txc_wr_pntr_1;
          txc_wr_pntr           <= txc_wr_pntr;
          compare_addr3_cmplt   <= '0';
        end if;
      end if;
    end if;
  end process;

-----------------------------------------------------------------------------
--  Generate address that will get the End Address
-----------------------------------------------------------------------------
  TXC_RD_ADDR : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if reset2tx_client = '1' then
        txc_mem_rd_addr       <= txc_min_rd_addr;
        txc_mem_rd_addr_0     <= txc_rd_addr5;
        txc_mem_rd_addr_1     <= txc_rd_addr6;
--  txc_rd_addr_cmp needs to lag one cnt because
--  it is incremented before the data is actually read
        txc_rd_addr_cmp       <= (others => '0');
      else
        if inc_txc_rd_addr = '1' and first_rd = '0' then
--  Initialize to start values
          txc_mem_rd_addr     <= txc_rd_addr5;
          txc_mem_rd_addr_0   <= txc_rd_addr6;
          txc_mem_rd_addr_1   <= txc_rd_addr7;
--  txc_rd_addr_cmp needs to lag one cnt because
--  it is incremented before the data is actually read
          txc_rd_addr_cmp     <= txc_min_rd_addr;
        elsif inc_txc_rd_addr = '1' and first_rd = '1' then
--  increment the address for the next packet
          if txc_mem_rd_addr = txc_max_rd_addr then
--  if the max address is reached, loop to address 0x4
            txc_mem_rd_addr   <= txc_mem_rd_addr_0;
            txc_mem_rd_addr_0 <= txc_mem_rd_addr_1;
            txc_mem_rd_addr_1 <= txc_rd_addr6;
            txc_rd_addr_cmp   <= txc_mem_rd_addr;
          else
--  otherwise just increment it
            txc_mem_rd_addr   <= txc_mem_rd_addr_0;
            txc_mem_rd_addr_0 <= txc_mem_rd_addr_1;
            txc_mem_rd_addr_1 <= std_logic_vector(unsigned(txc_mem_rd_addr_1) + 1);
            txc_rd_addr_cmp   <= txc_mem_rd_addr;
          end if;
        else                            -- Hold the current address until something changes
          txc_mem_rd_addr     <= txc_mem_rd_addr;
          txc_mem_rd_addr_0   <= txc_mem_rd_addr_0;
          txc_mem_rd_addr_1   <= txc_mem_rd_addr_1;
          txc_rd_addr_cmp     <= txc_rd_addr_cmp;
        end if;
      end if;
    end if;
  end process;


-----------------------------------------------------------------------------
--  Generate address mux fo memory
-----------------------------------------------------------------------------
  MEM_TXC_RD_ADDR : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if set_txc_addr4_n = '1' and first_rd = '0' and set_txc_wr = '0' then
-- Provide the address for the End of packet address
        Tx_Client_TxC_2_Mem_Addr_int <= txc_min_rd_addr;
      elsif set_txc_addr4_n = '1' and first_rd = '1' and set_txc_wr = '0' then
-- Provide the address for the End of packet address
        Tx_Client_TxC_2_Mem_Addr_int <= txc_mem_rd_addr;
      elsif set_txc_addr2 = '1' and set_txc_wr = '1' then
--Write the txc rd pointer
        Tx_Client_TxC_2_Mem_Addr_int <= txc_rd_addr2;
      elsif set_txc_addr3 = '1' and set_txc_wr = '0' then
--Read the txc wr pointer
        Tx_Client_TxC_2_Mem_Addr_int <= txc_rd_addr3;
      elsif set_txc_addr1 = '1' and set_txc_wr = '0' then
--  Read the TxD write pointer to monitor for an empty condition
        Tx_Client_TxC_2_Mem_Addr_int <= txc_rd_addr1;
      elsif set_txc_addr0 = '1' and set_txc_wr = '1' then
--  Write the current TxD Read Pointer while transmitting data
        Tx_Client_TxC_2_Mem_Addr_int <= txc_rd_addr0;
      else
        Tx_Client_TxC_2_Mem_Addr_int <= Tx_Client_TxC_2_Mem_Addr_int;
      end if;
    end if;
  end process;

  Tx_Client_TxC_2_Mem_Addr <= Tx_Client_TxC_2_Mem_Addr_int;

---------------------------------------------------------------------------
--  Write the TxC Rd Pointer to address 2 or
--    write the TxD Rd Pointer to address 0
--    Remove the lower 2 bits to align to a 32 bit word instead of a byte
---------------------------------------------------------------------------
  TXC_MEM_ADDR_PNTR : process(tx_axi_clk)
  begin
    if rising_edge(tx_axi_clk) then
      if set_txc_addr2 = '1' then
--Address for data that is currently being transmitted
        Tx_Client_TxC_2_Mem_Din_int <= zeroes_txc & txc_rd_addr_cmp(c_TxC_addra_width -1 downto 0);
      elsif set_txc_addr0 = '1' then
        Tx_Client_TxC_2_Mem_Din_int <= zeroes_txd & txd_rd_addr(c_TxD_addra_width -1 downto 2);
      else
        Tx_Client_TxC_2_Mem_Din_int <= (others => '0');
      end if;
    end if;
  end process;

  Tx_Client_TxC_2_Mem_Din <= Tx_Client_TxC_2_Mem_Din_int;

-----------------------------------------------------------------------------
--  Transmit Client TX Control State Machine Combinatorial Logic
-----------------------------------------------------------------------------
    FSM_TXCLIENT_TXD_CMB : process (txd_rd_cs,tx_axis_mac_tready,
        start_txd_fsm,
        Tx_Client_TxD_2_Mem_Dout, txd_rd_addr,txc_rd_end,
        end_addr, phy_mode_enable, enabled_1588,
        clr_txd_vld_d1)
    begin
        set_txd_vld      <= '0';
        clr_txd_vld      <= '0';
        set_txd_en       <= '0';
        inc_txd_rd_addr  <= '0';
        align_start_addr <= '0';
        set_txd_done     <= '0';
        load_tx_pipe     <= '0';
		flush_tx_pipe    <= '0';
        txd_rd_ns        <= txd_rd_cs;

        case txd_rd_cs is
            when IDLE       =>
                if start_txd_fsm = '1' then
                    set_txd_en      <= '1';
                    inc_txd_rd_addr <= '1';
                    txd_rd_ns       <= GET_B1;
                else
                    inc_txd_rd_addr <= '0';
                    set_txd_en      <= txc_rd_end;
                    txd_rd_ns       <= IDLE;
                end if;

            when GET_B1     =>
                inc_txd_rd_addr   <= '1';
                set_txd_vld       <= '1'; --Start sending first data of payload
                set_txd_en        <= '1';
                txd_rd_ns         <= STREAM_DATA;
            when WAIT_TRDY  =>
                if tx_axis_mac_tready = '1' then
	            flush_tx_pipe   <= '1';
		    if end_addr = txd_rd_addr then
                        if txd_rd_addr(1) = '1' and txd_rd_addr (0) = '1' then
                            align_start_addr <= '0';
                            inc_txd_rd_addr  <= '1';
                        else
                            align_start_addr <= '1';
                            inc_txd_rd_addr  <= '0';
                        end if;
                        if phy_mode_enable = '0' then
                            clr_txd_vld      <= '0';
                            set_txd_en       <= '0';
                            set_txd_done     <= '0';
                            txd_rd_ns        <= WAIT_LAST;
                        elsif phy_mode_enable = '1' then
                            clr_txd_vld      <= '1';
                            set_txd_en       <= '0';
                            set_txd_done     <= '1';
                            txd_rd_ns        <= IDLE;
                        end if;
                    else
                        inc_txd_rd_addr    <= '1'; 
                        set_txd_en         <= '1';
                        set_txd_done       <= '0';
                        align_start_addr   <= '0';
                        txd_rd_ns          <= STREAM_DATA;
                    end if;
                else
                    inc_txd_rd_addr <= '0';
                    set_txd_en      <= '0';
                    txd_rd_ns       <= WAIT_TRDY;
                end if;

            when STREAM_DATA =>
                if tx_axis_mac_tready = '1' then
--  The end addreess read from the memory is always one byte before
--  the actual end of the packet to allow tlast to be asserted correctly

--  On the write side of the BRAM, the end_addr has been set such that the
--  at strobes at TLAST reflect the last byte of data minus 1
--    case axi_str_txd_tstrb_dly0 is
--      when "1111" => end_addr_byte_offset <= "11";
--      when "0111" => end_addr_byte_offset <= "10";
--      when "0011" => end_addr_byte_offset <= "01";
--      when others => end_addr_byte_offset <= "00";
--    end case;
--
--  The BRAM parity bits are not used with AXI-S CORE Gen
--
                    if end_addr = txd_rd_addr then
--Last byte of payload data is one byte after end_address
                        if txd_rd_addr(1) = '1' and txd_rd_addr (0) = '1' then
--  By incrementing the address one, it will be 32 bit aligned
--  which is the starting address of the next packet
                            align_start_addr <= '0';
                            inc_txd_rd_addr  <= '1';
                        else
--  Align address to 32 bits because it ended non aligned
--    The next 32 bit aligned address will be the start
--    of the next payload data
--  Do not increment the address since it is getting aligned
                            align_start_addr <= '1';
                            inc_txd_rd_addr  <= '0';
                        end if;
                        if phy_mode_enable = '0' then
                            clr_txd_vld      <= '0';
                            set_txd_en       <= '0';
                            set_txd_done     <= '0';
                            txd_rd_ns        <= WAIT_LAST;
                        elsif phy_mode_enable = '1' then
                            clr_txd_vld      <= '1';
                            set_txd_en       <= '0';
                            set_txd_done     <= '1';
                            txd_rd_ns        <= IDLE;
                        end if;
                    else
                        inc_txd_rd_addr    <= '1'; --set addr to get next data
                        set_txd_en         <= '1';
                        set_txd_done       <= '0';
                        align_start_addr   <= '0';
                        txd_rd_ns          <= STREAM_DATA;
                    end if;
                else
                    inc_txd_rd_addr      <= '0';
                    set_txd_en           <= '0';
                    set_txd_done         <= '0';
                    align_start_addr     <= '0';
					load_tx_pipe         <= '1';
                    txd_rd_ns            <= WAIT_TRDY;
                end if;

            when WAIT_LAST =>
                if tx_axis_mac_tready = '1' and clr_txd_vld_d1 = '0' then
                    clr_txd_vld     <= '1';
                    inc_txd_rd_addr <= '0';
                    set_txd_en      <= '0';
                    set_txd_done    <= '0';
                    txd_rd_ns       <= WAIT_LAST;
		elsif tx_axis_mac_tready = '0' and clr_txd_vld_d1 = '0' then
                    clr_txd_vld     <= '0';
                    inc_txd_rd_addr <= '0';
                    set_txd_en      <= '0';
                    set_txd_done    <= '0';
                    txd_rd_ns       <= WAIT_LAST;
		elsif tx_axis_mac_tready = '1' and clr_txd_vld_d1 = '1' then	
				    clr_txd_vld     <= '0';
                    inc_txd_rd_addr <= '0';
                    set_txd_en      <= '0';
                    set_txd_done    <= '1';
                    txd_rd_ns       <= IDLE;
		elsif tx_axis_mac_tready = '1' and clr_txd_vld_d1 = '0' then	
				    clr_txd_vld     <= '1';
                    inc_txd_rd_addr <= '0';
                    set_txd_en      <= '0';
                    set_txd_done    <= '0';
                    txd_rd_ns       <= WAIT_LAST;	
                end if;    

            when others =>
                txd_rd_ns <= IDLE;

        end case;
    end process;

-----------------------------------------------------------------------------
--  Transmit Client TX Control State Machine Sequencer
-----------------------------------------------------------------------------
    FSM_TXCLIENT_TXD_SEQ : process (tx_axi_clk)
    begin
        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd_rd_cs <= IDLE;
            else
                txd_rd_cs <= txd_rd_ns;
            end if;
        end if;
    end process;


-----------------------------------------------------------------------------
--  Transmit Client TX Complete Signal
-----------------------------------------------------------------------------
    TX_COMPLETE_INDICATOR : process (tx_axi_clk)
    begin
        if rising_edge(tx_axi_clk) then
            if set_txd_done = '1' then
                tx_cmplt <= '1';
            else
                tx_cmplt <= '0';
            end if;
        end if;
    end process;


-----------------------------------------------------------------------------
--  Store 1 Byte in pipeline if tready is not asserted
-----------------------------------------------------------------------------
    TXD_BYTE1 : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd_pipe   <= (others => '0');
            else
                if load_tx_pipe = '1' then
                    txd_pipe <= Tx_Client_TxD_2_Mem_Dout(C_CLIENT_WIDTH-1 downto 0);
                else
                    txd_pipe <= txd_pipe;
                end if;
            end if;
        end if;
    end process;



-----------------------------------------------------------------------------
--  Use this delay to mux in the stored first bytes of data for each packet
-----------------------------------------------------------------------------
    TX_ACK_DELAY : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then

            if tx_axis_mac_tready = '1' then
                tx_axis_mac_tready_dly <= '1';
            else
                tx_axis_mac_tready_dly <= '0';
            end if;
        end if;

    end process;

-----------------------------------------------------------------------------
--  TxD Read Memory Enable - only enable memory when needed
-----------------------------------------------------------------------------
    TXD_MEM_EN : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if set_txd_en = '1' then
                Tx_Client_TxD_2_Mem_En_int <= '1';
            else
                Tx_Client_TxD_2_Mem_En_int <= '0';
            end if;
        end if;
    end process;

    Tx_Client_TxD_2_Mem_En <= Tx_Client_TxD_2_Mem_En_int;

-----------------------------------------------------------------------------
--  TxD Memory Write Enable bit is never written to
-----------------------------------------------------------------------------
    Tx_Client_TxD_2_Mem_We(0) <= '0';

-----------------------------------------------------------------------------
--  Get Lower 2 bits for case statement below
-----------------------------------------------------------------------------
    txd_rd_addr_1_0 <= txd_rd_addr(1 downto 0); -- for case statement below

-----------------------------------------------------------------------------
--  Set the address to be 32 bit aligned for readjustment at the end of
--    the packet
-----------------------------------------------------------------------------
  txd_rd_addr_aligned <= txd_rd_addr(c_TxD_addra_width -1 downto 2) & "00";

-----------------------------------------------------------------------------
--  Generate the TxD Memory Read Address
-----------------------------------------------------------------------------
      TXD_MEM_RD_ADDR : process(tx_axi_clk)
      begin
  
        if rising_edge(tx_axi_clk) then
          if reset2tx_client = '1' then
            txd_rd_addr     <= (others => '0');
          else
--  the end of the packet was reached, so adjust the Rd Addr
--    to be 32bit aligned if needed
            if align_start_addr = '1' then
              case txd_rd_addr_1_0 is
                when "00" | "01" | "10" => --  | "11" =>
-- packet ended on a non 32bit aligned address, so adjust it
                  txd_rd_addr <= std_logic_vector(unsigned(txd_rd_addr_aligned) + 4);
                when  others =>
-- packet ended on a 32bit aligned address, so do not change
                  txd_rd_addr <= txd_rd_addr;
              end case;
            else
--  increment to next address
              if inc_txd_rd_addr = '1' then
                txd_rd_addr <= std_logic_vector(unsigned(txd_rd_addr) + 1);
              else
                txd_rd_addr <= txd_rd_addr;
              end if;
            end if;
          end if;
        end if;
      end process;

        Tx_Client_TxD_2_Mem_Addr <= txd_rd_addr;


---------------------------------------------------------------------------
--  Force and update the BRAM with the rd_pntr_addr every ~512 bytes
---------------------------------------------------------------------------
    BRAM_UPDATE : process(tx_axi_clk)
    begin
        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' or set_txd_done = '1' then
                update_bram_cnt   <= (others => '0');
            else
                if update_bram_cnt(9) = '1' and inc_txd_rd_addr = '1' then
                    update_bram_cnt <= ('0' & update_bram_cnt(8 downto 0)) + 1;
                elsif inc_txd_rd_addr = '1' then
                    update_bram_cnt <= update_bram_cnt + 1;
                else
                    update_bram_cnt <= update_bram_cnt;
                end if;
            end if;
        end if;
    end process;


---------------------------------------------------------------------------
--  Use this signal to dis-allow a transition to the WAIT_TRDY3 state of
--  the FSM_TXCLIENT_TXD_CMB FSM when in the WAIT_TRDY2 state
---------------------------------------------------------------------------
        SET_FIRST_BYTE_FILTER : process (tx_axi_clk)
        begin
          if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
              clr_txd_vld_d1   <= '0';
            else
              if clr_txd_vld = '1' then
                clr_txd_vld_d1 <= '1';
			  else
                clr_txd_vld_d1 <= '0';
              end if;
            end if;
          end if;
        end process;


-----------------------------------------------------------------------------
--  Mux the Memory data to the Tx Client Interface when appropriate
--    1. Mux the first byte
--    2. Mux the second byte at the rising edge of the first tready of the packet
--    3. Mux the third byte at the second tready of the packet
--    4. Mux the fourth byte at the third tready of the packet
--    5. Mux the remaining bytes
-----------------------------------------------------------------------------
    TXD_MEM_DATA : process (tx_axi_clk)
    begin
        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd   <= (others => '0');
            else
                if set_txd_vld = '1' then
                    txd <= Tx_Client_TxD_2_Mem_Dout(C_CLIENT_WIDTH-1 downto 0); --load first byte and hold until ack
                elsif flush_tx_pipe = '1' then
				    txd <= txd_pipe; 
                elsif tx_axis_mac_tready = '1' then
                    txd <= Tx_Client_TxD_2_Mem_Dout(C_CLIENT_WIDTH -1 downto 0); --remaining bytes
                else
                    txd <= txd;
                end if;
            end if;
        end if;
    end process;

    tx_axis_mac_tdata <= txd;

-----------------------------------------------------------------------------
--  Assert Transmit Data Valid for the duration of a transmitted packet
-----------------------------------------------------------------------------
    SET_TX_DATA_VALID : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                txd_vld   <= '0';
            else
                if tx_axis_mac_tready = '1' and tx_axis_mac_tlast_int = '1' then
                    txd_vld <= '0';
                elsif set_txd_vld = '1' then
                    txd_vld <= '1';
                else
                    txd_vld <= txd_vld;
                end if;
            end if;
        end if;
    end process;

    tx_axis_mac_tvalid <= txd_vld;

-----------------------------------------------------------------------------
--  Assert Transmit Data LAST to end the packet
-----------------------------------------------------------------------------
    SET_TLAST : process (tx_axi_clk)
    begin

        if rising_edge(tx_axi_clk) then
            if reset2tx_client = '1' then
                tx_axis_mac_tlast_int   <= '0';
            elsif tx_axis_mac_tready = '1' then
                if clr_txd_vld = '1' then
                    tx_axis_mac_tlast_int <= '1';
                else
                    tx_axis_mac_tlast_int <= '0';
                end if;
            else
                tx_axis_mac_tlast_int   <= tx_axis_mac_tlast_int;
            end if;
        end if;
    end process;

    tx_axis_mac_tlast <= tx_axis_mac_tlast_int;


end rtl;


-------------------------------------------------------------------------------
-- tx_axistream_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_axistream_if.vhd
-- Version:         v1.00a
-- Description:     embedded ip AXI Stream transmit interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--          ->        tx_axistream_if.vhd
--                      tx_basic_if.vhd
--                      tx_csum_if.vhd
--                        tx_csum_partial_if.vhd
--                          tx_csum_partial_calc_if.vhd
--                        tx_full_csum_if.vhd
--                      tx_vlan_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd
--
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

library work;
use work.tx_if_pack.all;

-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity tx_axistream_if is
  generic (
    C_FAMILY               : string                       := "virtex6";
    C_HALFDUP              : integer range 0 to 1         := 0;
    C_TXCSUM               : integer range 0 to 2         := 0;
    C_TXMEM                : integer                      := 4096;
    C_TXVLAN_TRAN          : integer range 0 to 1         := 0;
    C_TXVLAN_TAG           : integer range 0 to 1         := 0;
    C_TXVLAN_STRP          : integer range 0 to 1         := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32       := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32       := 32;

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    : integer range  36 to 36     := 36;
    c_TxD_read_width_b     : integer range  36 to 36     := 36;
    c_TxD_write_depth_b    : integer range   0 to 8192   := 4096;
    c_TxD_read_depth_b     : integer range   0 to 8192   := 4096;
    c_TxD_addrb_width      : integer range   0 to 13     := 10;
    c_TxD_web_width        : integer range   0 to 4      := 4;

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    : integer range   36 to 36    := 36;
    c_TxC_read_width_b     : integer range   36 to 36    := 36;
    c_TxC_write_depth_b    : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b     : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width      : integer range    0 to 10    := 10;
    c_TxC_web_width        : integer range    0 to 1     := 1
  );
  port (

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       : in  std_logic;                                           --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      : in  std_logic;                                           --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     : in  std_logic;                                           --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     : out std_logic;                                           --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      : in  std_logic;                                           --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      : in  std_logic_vector(3 downto 0);                        --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);     --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       : in  std_logic;                                           --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      : in  std_logic;                                           --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     : in  std_logic;                                           --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     : out std_logic;                                           --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      : in  std_logic;                                           --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      : in  std_logic_vector(3 downto 0);                        --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);     --  AXI-Stream Transmit Control Data


    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  : out std_logic_vector(c_TxD_write_width_b-1 downto 0);    --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr : out std_logic_vector(c_TxD_addrb_width-1   downto 0);    --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   : out std_logic;                                           --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   : out std_logic_vector(c_TxD_web_width-1     downto 0);    --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout : in  std_logic_vector(c_TxD_read_width_b-1  downto 0);    --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  : out std_logic_vector(c_TxC_write_width_b-1 downto 0);    --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr : out std_logic_vector(c_TxC_addrb_width-1   downto 0);    --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   : out std_logic;                                           --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   : out std_logic_vector(c_TxC_web_width-1     downto 0);    --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout : in  std_logic_vector(c_TxC_read_width_b-1  downto 0);    --  Tx AXI-Stream Control to Memory Full Flag

    -- VLAN Signals
    tx_vlan_bram_addr      : out std_logic_vector(11 downto 0);                       --  Transmit VLAN BRAM Addr
    tx_vlan_bram_din       : in  std_logic_vector(13 downto 0);                       --  Transmit VLAN BRAM Rd Data
    tx_vlan_bram_en        : out std_logic;                                           --  Transmit VLAN BRAM Enable

    enable_newFncEn        : out std_logic; --Only perform VLAN when the FLAG = 0xA   --  Enable Extended VLAN Functions
    transMode_cross        : in  std_logic;                                           --  VLAN Translation Mode Control Bit
    tagMode_cross          : in  std_logic_vector( 1 downto 0);                       --  VLAN TAG Mode Control Bits
    strpMode_cross         : in  std_logic_vector( 1 downto 0);                       --  VLAN Strip Mode Control Bits

    tpid0_cross            : in  std_logic_vector(15 downto 0);                       --  VLAN TPID
    tpid1_cross            : in  std_logic_vector(15 downto 0);                       --  VLAN TPID
    tpid2_cross            : in  std_logic_vector(15 downto 0);                       --  VLAN TPID
    tpid3_cross            : in  std_logic_vector(15 downto 0);                       --  VLAN TPID

    newTagData_cross       : in  std_logic_vector(31 downto 0);                       --  VLAN Tag Data

    tx_init_in_prog        : out std_logic                                            --  Tx is Initializing after a reset

  );

end tx_axistream_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of tx_axistream_if is

begin

-------------------------------------------------------------------------------
--  Start Basic Design - No CSUM,  No Extended VLAN
-------------------------------------------------------------------------------
GEN_BASIC : if ( (C_TXCSUM  = 0 and (C_TXVLAN_TRAN = 0 and C_TXVLAN_TAG = 0 and C_TXVLAN_STRP = 0)) or
                 (C_TXCSUM /= 0 and (C_TXVLAN_TRAN = 1  or C_TXVLAN_TAG = 1  or C_TXVLAN_STRP = 1))) generate
begin


  tx_vlan_bram_addr <= (others => '0');
  tx_vlan_bram_en   <= '0';
  enable_newFncEn   <= '0';

  TX_BASIC_INTERFACE : tx_basic_if
  --  Interface for Transmit AxiStream Data and Control; and Tx Memory
  generic map (
    C_FAMILY               => C_FAMILY,
    C_HALFDUP              => C_HALFDUP,
    C_TXCSUM               => C_TXCSUM,
    C_TXMEM                => C_TXMEM,
    C_TXVLAN_TRAN          => C_TXVLAN_TRAN,
    C_TXVLAN_TAG           => C_TXVLAN_TAG,
    C_TXVLAN_STRP          => C_TXVLAN_STRP,
    C_S_AXI_ADDR_WIDTH     => C_S_AXI_ADDR_WIDTH,
    C_S_AXI_DATA_WIDTH     => C_S_AXI_DATA_WIDTH,

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    => c_TxD_write_width_b,
    c_TxD_read_width_b     => c_TxD_read_width_b,
    c_TxD_write_depth_b    => c_TxD_write_depth_b,
    c_TxD_read_depth_b     => c_TxD_read_depth_b,
    c_TxD_addrb_width      => c_TxD_addrb_width,
    c_TxD_web_width        => c_TxD_web_width,

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    => c_TxC_write_width_b,
    c_TxC_read_width_b     => c_TxC_read_width_b,
    c_TxC_write_depth_b    => c_TxC_write_depth_b,
    c_TxC_read_depth_b     => c_TxC_read_depth_b,
    c_TxC_addrb_width      => c_TxC_addrb_width,
    c_TxC_web_width        => c_TxC_web_width

  )
  port map  (

    tx_init_in_prog        => tx_init_in_prog,             --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       => AXI_STR_TXD_ACLK,            --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      => reset2axi_str_txd,           --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     => AXI_STR_TXD_TVALID,          --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     => AXI_STR_TXD_TREADY,          --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      => AXI_STR_TXD_TLAST,           --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      => AXI_STR_TXD_TSTRB,           --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      => AXI_STR_TXD_TDATA,           --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       => AXI_STR_TXC_ACLK,            --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      => reset2axi_str_txc,           --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     => AXI_STR_TXC_TVALID,          --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     => AXI_STR_TXC_TREADY,          --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      => AXI_STR_TXC_TLAST,           --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      => AXI_STR_TXC_TSTRB,           --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      => AXI_STR_TXC_TDATA,           --  AXI-Stream Transmit Control Data

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  => Axi_Str_TxD_2_Mem_Din,       --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr => Axi_Str_TxD_2_Mem_Addr,      --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   => Axi_Str_TxD_2_Mem_En,        --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   => Axi_Str_TxD_2_Mem_We,        --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout => Axi_Str_TxD_2_Mem_Dout,      --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  => Axi_Str_TxC_2_Mem_Din,       --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr => Axi_Str_TxC_2_Mem_Addr,      --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   => Axi_Str_TxC_2_Mem_En,        --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   => Axi_Str_TxC_2_Mem_We,        --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout => Axi_Str_TxC_2_Mem_Dout       --  Tx AXI-Stream Control to Memory Full Flag

  );

end generate GEN_BASIC;
-------------------------------------------------------------------------------
--  End Basic Design
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
--  Start CSUM
-------------------------------------------------------------------------------
GEN_CSUM : if (C_TXCSUM  = 1 and (C_TXVLAN_TRAN = 0 and C_TXVLAN_TAG = 0 and C_TXVLAN_STRP = 0)) or
              (C_TXCSUM  = 2 and (C_TXVLAN_TRAN = 0 and C_TXVLAN_TAG = 0 and C_TXVLAN_STRP = 0)) generate
begin


  tx_vlan_bram_addr <= (others => '0');
  tx_vlan_bram_en   <= '0';
  enable_newFncEn   <= '0';

  TX_CSUM_INTERFACE : tx_csum_if
  --  Interface for Transmit AxiStream Data and Control; and Tx Memory
  generic map (
    C_FAMILY               => C_FAMILY,
    C_HALFDUP              => C_HALFDUP,
    C_TXCSUM               => C_TXCSUM,
    C_TXMEM                => C_TXMEM,
    C_TXVLAN_TRAN          => C_TXVLAN_TRAN,
    C_TXVLAN_TAG           => C_TXVLAN_TAG,
    C_TXVLAN_STRP          => C_TXVLAN_STRP,
    C_S_AXI_ADDR_WIDTH     => C_S_AXI_ADDR_WIDTH,
    C_S_AXI_DATA_WIDTH     => C_S_AXI_DATA_WIDTH,

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    => c_TxD_write_width_b,
    c_TxD_read_width_b     => c_TxD_read_width_b,
    c_TxD_write_depth_b    => c_TxD_write_depth_b,
    c_TxD_read_depth_b     => c_TxD_read_depth_b,
    c_TxD_addrb_width      => c_TxD_addrb_width,
    c_TxD_web_width        => c_TxD_web_width,

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    => c_TxC_write_width_b,
    c_TxC_read_width_b     => c_TxC_read_width_b,
    c_TxC_write_depth_b    => c_TxC_write_depth_b,
    c_TxC_read_depth_b     => c_TxC_read_depth_b,
    c_TxC_addrb_width      => c_TxC_addrb_width,
    c_TxC_web_width        => c_TxC_web_width

  )
  port map  (

    tx_init_in_prog        => tx_init_in_prog,             --  Tx is Initializing after a reset

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK       => AXI_STR_TXD_ACLK,            --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd      => reset2axi_str_txd,           --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID     => AXI_STR_TXD_TVALID,          --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY     => AXI_STR_TXD_TREADY,          --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST      => AXI_STR_TXD_TLAST,           --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB      => AXI_STR_TXD_TSTRB,           --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA      => AXI_STR_TXD_TDATA,           --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       => AXI_STR_TXC_ACLK,            --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      => reset2axi_str_txc,           --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     => AXI_STR_TXC_TVALID,          --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     => AXI_STR_TXC_TREADY,          --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      => AXI_STR_TXC_TLAST,           --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      => AXI_STR_TXC_TSTRB,           --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      => AXI_STR_TXC_TDATA,           --  AXI-Stream Transmit Control Data

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  => Axi_Str_TxD_2_Mem_Din,
    Axi_Str_TxD_2_Mem_Addr => Axi_Str_TxD_2_Mem_Addr,      --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_En   => Axi_Str_TxD_2_Mem_En,        --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_We   => Axi_Str_TxD_2_Mem_We,        --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_Dout => Axi_Str_TxD_2_Mem_Dout,      --  Tx AXI-Stream Data to Memory Wr En
                                                           --  Tx AXI-Stream Data to Memory Not Used
    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  => Axi_Str_TxC_2_Mem_Din,
    Axi_Str_TxC_2_Mem_Addr => Axi_Str_TxC_2_Mem_Addr,      --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_En   => Axi_Str_TxC_2_Mem_En,        --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_We   => Axi_Str_TxC_2_Mem_We,        --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_Dout => Axi_Str_TxC_2_Mem_Dout       --  Tx AXI-Stream Control to Memory Wr En
                                                           --  Tx AXI-Stream Control to Memory Full Flag
  );

end generate GEN_CSUM;
-------------------------------------------------------------------------------
--  End CSUM
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
--  Start Extended VLAN
-------------------------------------------------------------------------------
GEN_EXT_VLAN : if ( C_TXCSUM  = 0 and (C_TXVLAN_TRAN = 1 or C_TXVLAN_TAG = 1 or C_TXVLAN_STRP = 1)) generate
begin

  TX_VLAN_INTERFACE : tx_vlan_if
  generic map (
    C_FAMILY               => C_FAMILY,
    C_HALFDUP              => C_HALFDUP,
    C_TXCSUM               => C_TXCSUM,
    C_TXMEM                => C_TXMEM,
    C_TXVLAN_TRAN          => C_TXVLAN_TRAN,
    C_TXVLAN_TAG           => C_TXVLAN_TAG,
    C_TXVLAN_STRP          => C_TXVLAN_STRP,
    C_S_AXI_ADDR_WIDTH     => C_S_AXI_ADDR_WIDTH,
    C_S_AXI_DATA_WIDTH     => C_S_AXI_DATA_WIDTH,

    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b    => c_TxD_write_width_b,
    c_TxD_read_width_b     => c_TxD_read_width_b,
    c_TxD_write_depth_b    => c_TxD_write_depth_b,
    c_TxD_read_depth_b     => c_TxD_read_depth_b,
    c_TxD_addrb_width      => c_TxD_addrb_width,
    c_TxD_web_width        => c_TxD_web_width,

    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b    => c_TxC_write_width_b,
    c_TxC_read_width_b     => c_TxC_read_width_b,
    c_TxC_write_depth_b    => c_TxC_write_depth_b,
    c_TxC_read_depth_b     => c_TxC_read_depth_b,
    c_TxC_addrb_width      => c_TxC_addrb_width,
    c_TxC_web_width        => c_TxC_web_width

  )
  port map  (

    tx_init_in_prog        => tx_init_in_prog,        --  Tx is Initializing after a reset

    -- AXI Stream Data signals                        --  AXI-Stream Transmit Data Clk
    AXI_STR_TXD_ACLK       => AXI_STR_TXD_ACLK,       --  AXI-Stream Transmit Data Reset
    reset2axi_str_txd      => reset2axi_str_txd,      --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TVALID     => AXI_STR_TXD_TVALID,     --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TREADY     => AXI_STR_TXD_TREADY,     --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TLAST      => AXI_STR_TXD_TLAST,      --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TSTRB      => AXI_STR_TXD_TSTRB,      --  AXI-Stream Transmit Data Data
    AXI_STR_TXD_TDATA      => AXI_STR_TXD_TDATA,
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK       => AXI_STR_TXC_ACLK,       --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc      => reset2axi_str_txc,      --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID     => AXI_STR_TXC_TVALID,     --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY     => AXI_STR_TXC_TREADY,     --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST      => AXI_STR_TXC_TLAST,      --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB      => AXI_STR_TXC_TSTRB,      --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA      => AXI_STR_TXC_TDATA,      --  AXI-Stream Transmit Control Data

    -- Write Port - AXI Stream TxData
    Axi_Str_TxD_2_Mem_Din  => Axi_Str_TxD_2_Mem_Din,  --  Tx AXI-Stream Data to Memory Wr Din
    Axi_Str_TxD_2_Mem_Addr => Axi_Str_TxD_2_Mem_Addr, --  Tx AXI-Stream Data to Memory Wr Addr
    Axi_Str_TxD_2_Mem_En   => Axi_Str_TxD_2_Mem_En,   --  Tx AXI-Stream Data to Memory Enable
    Axi_Str_TxD_2_Mem_We   => Axi_Str_TxD_2_Mem_We,   --  Tx AXI-Stream Data to Memory Wr En
    Axi_Str_TxD_2_Mem_Dout => Axi_Str_TxD_2_Mem_Dout, --  Tx AXI-Stream Data to Memory Not Used

    -- Write Port - AXI Stream TxControl
    Axi_Str_TxC_2_Mem_Din  => Axi_Str_TxC_2_Mem_Din,  --  Tx AXI-Stream Control to Memory Wr Din
    Axi_Str_TxC_2_Mem_Addr => Axi_Str_TxC_2_Mem_Addr, --  Tx AXI-Stream Control to Memory Wr Addr
    Axi_Str_TxC_2_Mem_En   => Axi_Str_TxC_2_Mem_En,   --  Tx AXI-Stream Control to Memory Enable
    Axi_Str_TxC_2_Mem_We   => Axi_Str_TxC_2_Mem_We,   --  Tx AXI-Stream Control to Memory Wr En
    Axi_Str_TxC_2_Mem_Dout => Axi_Str_TxC_2_Mem_Dout, --  Tx AXI-Stream Control to Memory Full Flag

    tx_vlan_bram_addr      => tx_vlan_bram_addr,      --  Transmit VLAN BRAM Addr
    tx_vlan_bram_din       => tx_vlan_bram_din,       --  Transmit VLAN BRAM Rd Data
    tx_vlan_bram_en        => tx_vlan_bram_en,        --  Transmit VLAN BRAM Enable

    enable_newFncEn        => enable_newFncEn,        --  Enable Extended VLAN Functions
    transMode_cross        => transMode_cross,        --  VLAN Translation Mode Control Bit
    tagMode_cross          => tagMode_cross,          --  VLAN TAG Mode Control Bits
    strpMode_cross         => strpMode_cross,         --  VLAN Strip Mode Control Bits

    tpid0_cross            => tpid0_cross,            --  VLAN TPID
    tpid1_cross            => tpid1_cross,            --  VLAN TPID
    tpid2_cross            => tpid2_cross,            --  VLAN TPID
    tpid3_cross            => tpid3_cross,            --  VLAN TPID

    newTagData_cross       => newTagData_cross        --  VLAN Tag Data
    );

end generate GEN_EXT_VLAN;
-------------------------------------------------------------------------------
--  Start Extended VLAN
-------------------------------------------------------------------------------
end rtl;


------------------------------------------------------------------------------
-- addr_response_shim.vhd
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        addr_response_shim.vhd
-- Version:         v1.00a
-- Description:     address response shim
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--            -- xps_ll_temac.vhd
--               -- addr_response_shim.vhd    ******
--               -- axi_soft_temac_wrap.vhd
--               -- v6_temac_wrap.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.

------------------------------------------------------------------------------
-- Author:
-- History:
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.all;

-------------------------------------------------------------------------------
-- Entity section
-------------------------------------------------------------------------------

entity addr_response_shim is
   generic (

      C_BUS2CORE_CLK_RATIO      : integer range 1 to 2    := 1;
      C_S_AXI_ADDR_WIDTH        : integer range 32 to 32  := 32;
      C_S_AXI_DATA_WIDTH        : integer range 32 to 32  := 32;
      C_SIPIF_DWIDTH            : integer range 32 to 32  := 32;
      C_NUM_CS                  : integer                 := 10;
      C_NUM_CE                  : integer                 := 41;
      C_FAMILY                  : string                  := "virtex6"
      );
   port (
      --Clock and Reset
      BUS2IP_CLK                : in  std_logic;                                        --  AXI4-Lite clk
      BUS2IP_RESET              : in  std_logic;                                        --  AXI4-Lite reset

      -- PLB Slave Interface with Shim
      BUS2IP_Addr               : in  std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );   --  Address bus from AXI4-Lite to Shim
      BUS2IP_Data               : in  std_logic_vector(0 to C_SIPIF_DWIDTH - 1 );       --  Data bus from AXI4-Lite to Shim
      BUS2IP_RNW                : in  std_logic;                                        --  RNW signal from AXI4-Lite to Shim
      BUS2IP_CS                 : in  std_logic_vector(0 to 0);                         --  CS signal from AXI4-Lite to Shim
      BUS2IP_RdCE               : in  std_logic_vector(0 to 0);                         --  RdCE signal from AXI4-Lite to Shim
      BUS2IP_WrCE               : in  std_logic_vector(0 to 0);                         --  WrCE signal from AXI4-Lite to Shim

      IP2BUS_Data               : out std_logic_vector (0 to C_SIPIF_DWIDTH - 1 );      --  Data bus from Shim to AXI4-Lite
      IP2BUS_WrAck              : out std_logic;                                        --  WrCE signal from Shim to AXI4-Lite
      IP2BUS_RdAck              : out std_logic;                                        --  RdCE signal from Shim to AXI4-Lite

      -- TEMAC Interface with Shim
      Shim2IP_Addr              : out std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );   --  Address bus from Shim to AXI Ethernet
      Shim2IP_Data              : out std_logic_vector(0 to C_SIPIF_DWIDTH - 1 );       --  Data bus from Shim to AXI Ethernet
      Shim2IP_RNW               : out std_logic;                                        --  RNW signal from Shim to AXI Ethernet
      Shim2IP_CS                : out std_logic_vector(0 to C_NUM_CS);                  --  CS signal from Shim to AXI Ethernet
      Shim2IP_RdCE              : out std_logic_vector(0 to C_NUM_CE);                  --  RdCE signal from Shim to AXI Ethernet
      Shim2IP_WrCE              : out std_logic_vector(0 to C_NUM_CE);                  --  WrCE signal from Shim to AXI Ethernet

      IP2Shim_Data              : in  std_logic_vector (0 to C_SIPIF_DWIDTH - 1 );      --  Data bus from AXI Ethernet to Shim
      IP2Shim_WrAck             : in  std_logic;                                        --  WrCE signal from AXI Ethernet to Shim
      IP2Shim_RdAck             : in  std_logic                                         --  RdCE signal from AXI Ethernet to Shim
   );

end addr_response_shim;

architecture rtl of addr_response_shim is


   signal BUS2IP_Addr_reg    : std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );
   signal BUS2IP_CS_reg      : std_logic;
   signal shim2IP_RNW_int      : std_logic;
   signal BUS2IP_RdCE_reg    : std_logic;
   signal BUS2IP_WrCE_reg    : std_logic;
   signal invalidAddrRspns     : std_logic;
   signal invalidAddrRspns_reg : std_logic;
   signal invalidRdReq         : std_logic;
   signal invalidWrReq         : std_logic;
   signal shim2IP_CS_int       : std_logic_vector(0 to C_NUM_CS);
   signal shim2IP_RdCE_int     : std_logic_vector(0 to C_NUM_CE);
   signal shim2IP_WrCE_int     : std_logic_vector(0 to C_NUM_CE);
   signal IP2Shim_WrAck_int    : std_logic;
   signal IP2Shim_RdAck_int    : std_logic;

   begin


      IP2Shim_WrAck_int <= IP2Shim_WrAck or invalidWrReq;
      IP2Shim_RdAck_int <= IP2Shim_RdAck or invalidRdReq;

      Shim2IP_Data      <= BUS2IP_Data ;  --write data

      IP2BUS_Data     <= IP2Shim_Data;    --read data
      IP2BUS_WrAck    <= IP2Shim_WrAck_int;
      IP2BUS_RdAck    <= IP2Shim_rDAck_int;

      ----------------------------------------------------------------------------
      -- Use Chip Select to register the address data; Otherwise Zeros
      ----------------------------------------------------------------------------
      ADDR_REG : process (BUS2IP_CLK)
      begin

         if rising_edge(BUS2IP_CLK) then
            if BUS2IP_RESET = '1' or (IP2Shim_WrAck_int = '1' or IP2Shim_RdAck_int = '1') then
               BUS2IP_Addr_reg <= (others => '0');
            elsif BUS2IP_CS(0) = '1' then
               BUS2IP_Addr_reg <= BUS2IP_Addr;
            else
               BUS2IP_Addr_reg <= BUS2IP_Addr_reg;
            end if;
         end if;
      end process;

      ----------------------------------------------------------------------------
      -- Use Chip Select to register Chip Select; Otherwise Zero
      ----------------------------------------------------------------------------
      CS_REG : process (BUS2IP_CLK)
      begin

         if rising_edge(BUS2IP_CLK) then
            if BUS2IP_RESET = '1' or (IP2Shim_WrAck_int = '1' or IP2Shim_RdAck_int = '1') then
               BUS2IP_CS_reg <= '0';
            elsif BUS2IP_CS(0) = '1' then
               BUS2IP_CS_reg <= BUS2IP_CS(0);
            else
               BUS2IP_CS_reg <= BUS2IP_CS_reg;
            end if;
         end if;
      end process;

      ----------------------------------------------------------------------------
      -- Use Chip Select to register Read Not Write; Otherwise Zero
      ----------------------------------------------------------------------------
      RNW_REG : process (BUS2IP_CLK)
      begin

         if rising_edge(BUS2IP_CLK) then
            if BUS2IP_RESET = '1' or (IP2Shim_WrAck_int = '1' or IP2Shim_RdAck_int = '1') then
               shim2IP_RNW_int <= '0';
            elsif BUS2IP_CS(0) = '1' then
               shim2IP_RNW_int <= BUS2IP_RNW;
            else
               shim2IP_RNW_int <= shim2IP_RNW_int;
            end if;
         end if;
      end process;

      ----------------------------------------------------------------------------
      -- Use Chip Select and BUS2IP_RNW to register Read Chip Enable
      -- Otherwise Zero
      ----------------------------------------------------------------------------
      RDCE_REG : process (BUS2IP_CLK)
      begin

         if rising_edge(BUS2IP_CLK) then
            if BUS2IP_RESET = '1' or (IP2Shim_WrAck_int = '1' or IP2Shim_RdAck_int = '1') then
               BUS2IP_RdCE_reg <= '0';
            elsif BUS2IP_CS(0) = '1' and BUS2IP_RNW = '1' then
               BUS2IP_RdCE_reg <= BUS2IP_RdCE(0);
            else
               BUS2IP_RdCE_reg <= BUS2IP_RdCE_reg;
            end if;
         end if;
      end process;

      ----------------------------------------------------------------------------
      -- Use Chip Select and BUS2IP_RNW to register Write Chip Enable
      -- Otherwise Zero
      ----------------------------------------------------------------------------
      WRCE_REG : process (BUS2IP_CLK)
      begin

         if rising_edge(BUS2IP_CLK) then
            if BUS2IP_RESET = '1' or (IP2Shim_WrAck_int = '1' or IP2Shim_RdAck_int = '1') then
               BUS2IP_WrCE_reg <= '0';
            elsif BUS2IP_CS(0) = '1' and BUS2IP_RNW = '0' then
               BUS2IP_WrCE_reg <= BUS2IP_WrCE(0);
            else
               BUS2IP_WrCE_reg <= BUS2IP_WrCE_reg;
            end if;
         end if;
      end process;


      ----------------------------------------------------------------------------
      -- Decode the address and set appropriate CE
      --    If the Address does not exist, ie it is in a gap,
      --    then set invalidAddrRspns
      ----------------------------------------------------------------------------
      ADDR_DECODE : process (BUS2IP_CS_reg,BUS2IP_RdCE_reg,BUS2IP_WrCE_reg,
                             BUS2IP_Addr_reg)
      begin


         if BUS2IP_CS_reg = '1' then
            if BUS2IP_Addr_reg(14 to 29) = "0000000000000000" then   --0x0
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- RAF
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(0)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(1 to C_NUM_CE)   <= (others => '0');
               shim2IP_WrCE_int(1 to C_NUM_CE)   <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000000001" then --0x4
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- TPF
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0)               <= '0';
               shim2IP_WrCE_int(0)               <= '0';
               shim2IP_RdCE_int(1)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(1)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(2 to C_NUM_CE)   <= (others => '0');
               shim2IP_WrCE_int(2 to C_NUM_CE)   <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000000010" then --0x8
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- IFGP
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 1)          <= (others => '0');
               shim2IP_WrCE_int(0 to 1)          <= (others => '0');
               shim2IP_RdCE_int(2)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(2)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(3 to C_NUM_CE)   <= (others => '0');
               shim2IP_WrCE_int(3 to C_NUM_CE)   <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000000011" then --0xC
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- IS
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 2)          <= (others => '0');
               shim2IP_WrCE_int(0 to 2)          <= (others => '0');
               shim2IP_RdCE_int(3)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(3)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(4 to C_NUM_CE)   <= (others => '0');
               shim2IP_WrCE_int(4 to C_NUM_CE)   <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000000100" then --0x10
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- IP
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 3)          <= (others => '0');
               shim2IP_WrCE_int(0 to 3)          <= (others => '0');
               shim2IP_RdCE_int(4)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(4)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(5 to C_NUM_CE)   <= (others => '0');
               shim2IP_WrCE_int(5 to C_NUM_CE)   <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000000101" then --0x14
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- IE
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 4)          <= (others => '0');
               shim2IP_WrCE_int(0 to 4)          <= (others => '0');
               shim2IP_RdCE_int(5)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(5)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(6 to C_NUM_CE)   <= (others => '0');
               shim2IP_WrCE_int(6 to C_NUM_CE)   <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000000110" then --0x18
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- TTAG
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 5)          <= (others => '0');
               shim2IP_WrCE_int(0 to 5)          <= (others => '0');
               shim2IP_RdCE_int(6)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(6)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(7 to C_NUM_CE)   <= (others => '0');
               shim2IP_WrCE_int(7 to C_NUM_CE)   <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000000111" then --0x1C
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- RTAG
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 6)          <= (others => '0');
               shim2IP_WrCE_int(0 to 6)          <= (others => '0');
               shim2IP_RdCE_int(7)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(7)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(8 to C_NUM_CE)   <= (others => '0');
               shim2IP_WrCE_int(8 to C_NUM_CE)   <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000001000" then --0x20
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- UAWL
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 7)          <= (others => '0');
               shim2IP_WrCE_int(0 to 7)          <= (others => '0');
               shim2IP_RdCE_int(8)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(8)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(9 to C_NUM_CE)   <= (others => '0');
               shim2IP_WrCE_int(9 to C_NUM_CE)   <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000001001" then --0x24
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- UAWU
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 8)          <= (others => '0');
               shim2IP_WrCE_int(0 to 8)          <= (others => '0');
               shim2IP_RdCE_int(9)               <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(9)               <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(10 to C_NUM_CE)  <= (others => '0');
               shim2IP_WrCE_int(10 to C_NUM_CE)  <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000001010" then --0x28
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- TPID0
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 9)          <= (others => '0');
               shim2IP_WrCE_int(0 to 9)          <= (others => '0');
               shim2IP_RdCE_int(10)              <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(10)              <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(11 to C_NUM_CE)  <= (others => '0');
               shim2IP_WrCE_int(11 to C_NUM_CE)  <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000001011" then --0x2C
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- TPID1
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 10)         <= (others => '0');
               shim2IP_WrCE_int(0 to 10)         <= (others => '0');
               shim2IP_RdCE_int(11)              <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(11)              <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(12 to C_NUM_CE)  <= (others => '0');
               shim2IP_WrCE_int(12 to C_NUM_CE)  <= (others => '0');
               invalidAddrRspns                  <= '0';
            elsif BUS2IP_Addr_reg(14 to 29) = "0000000000001100" then --0x30
               shim2IP_CS_int(0)                 <= BUS2IP_CS_reg;      -- PCSPMA Status
               shim2IP_CS_int(1 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 11)         <= (others => '0');
               shim2IP_WrCE_int(0 to 11)         <= (others => '0');
               shim2IP_RdCE_int(12)              <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(12)              <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(13 to C_NUM_CE)  <= (others => '0');
               shim2IP_WrCE_int(13 to C_NUM_CE)  <= (others => '0');
               invalidAddrRspns                  <= '0';

            -- statistics and temac registers via external shim decode
            elsif BUS2IP_Addr_reg(14 to 22) = "000000001" or
                  BUS2IP_Addr_reg(14 to 21) = "00000001" then        --0x00200 - 0x007FC
               shim2IP_CS_int(0)                 <= '0';
               shim2IP_CS_int(1)                 <= BUS2IP_CS_reg;
               shim2IP_CS_int(2 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 15)         <= (others => '0');
               shim2IP_WrCE_int(0 to 15)         <= (others => '0');
               shim2IP_RdCE_int(16)              <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(16)              <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(17 to C_NUM_CE)  <= (others => '0');
               shim2IP_WrCE_int(17 to C_NUM_CE)  <= (others => '0');
               invalidAddrRspns                  <= '0';
            -- Tx VLAN
            elsif BUS2IP_Addr_reg(14 to 17) = "0001" then        --0x04000 - 0x07FFC
               shim2IP_CS_int(0 to 1)            <= (others => '0');
               shim2IP_CS_int(2)                 <= BUS2IP_CS_reg;
               shim2IP_CS_int(3 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 16)         <= (others => '0');
               shim2IP_WrCE_int(0 to 16)         <= (others => '0');
               shim2IP_RdCE_int(17)              <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(17)              <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(18 to C_NUM_CE)  <= (others => '0');
               shim2IP_WrCE_int(18 to C_NUM_CE)  <= (others => '0');
               invalidAddrRspns                  <= '0';
            -- Rx VLAN
            elsif BUS2IP_Addr_reg(14 to 16) = "001" then        --0x08000 - 0x0BFFC
               shim2IP_CS_int(0 to 2)            <= (others => '0');
               shim2IP_CS_int(3)                 <= BUS2IP_CS_reg;
               shim2IP_CS_int(4 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 17)         <= (others => '0');
               shim2IP_WrCE_int(0 to 17)         <= (others => '0');
               shim2IP_RdCE_int(18)              <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(18)              <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(19 to C_NUM_CE)  <= (others => '0');
               shim2IP_WrCE_int(19 to C_NUM_CE)  <= (others => '0');
               invalidAddrRspns                  <= '0';
            -- AVB
            elsif BUS2IP_Addr_reg(14 to 15) = "01" then        --0x010000 - 0x013FFC
               shim2IP_CS_int(0 to 3)            <= (others => '0');
               shim2IP_CS_int(4)                 <= BUS2IP_CS_reg;
               shim2IP_CS_int(5 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 18)         <= (others => '0');
               shim2IP_WrCE_int(0 to 18)         <= (others => '0');
               shim2IP_RdCE_int(19)              <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(19)              <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(20 to C_NUM_CE)  <= (others => '0');
               shim2IP_WrCE_int(20 to C_NUM_CE)  <= (others => '0');
               invalidAddrRspns                  <= '0';
            -- multicast
            elsif BUS2IP_Addr_reg(14) = '1' then        --0x020000 - 0x03FFFC
               shim2IP_CS_int(0 to 4)            <= (others => '0');
               shim2IP_CS_int(5)                 <= BUS2IP_CS_reg;
               shim2IP_CS_int(6 to C_NUM_CS)     <= (others => '0');
               shim2IP_RdCE_int(0 to 19)         <= (others => '0');
               shim2IP_WrCE_int(0 to 19)         <= (others => '0');
               shim2IP_RdCE_int(20)              <= BUS2IP_RdCE_reg;
               shim2IP_WrCE_int(20)              <= BUS2IP_WrCE_reg;
               shim2IP_RdCE_int(21 to C_NUM_CE)  <= (others => '0');
               shim2IP_WrCE_int(21 to C_NUM_CE)  <= (others => '0');
               invalidAddrRspns                  <= '0';
            else
               shim2IP_CS_int       <= (others => '0');
               shim2IP_RdCE_int     <= (others => '0');
               shim2IP_WrCE_int     <= (others => '0');
               invalidAddrRspns     <= '1';
            end if;
         else
            shim2IP_CS_int       <= (others => '0');
            shim2IP_RdCE_int     <= (others => '0');
            shim2IP_WrCE_int     <= (others => '0');
            invalidAddrRspns     <= '0';
         end if;
      end process;


      ----------------------------------------------------------------------------
      -- Register Address Decode Signals for timing
      ----------------------------------------------------------------------------
      REG_DECODE_SIGNALS : process (BUS2IP_CLK)
      begin

         if rising_edge(BUS2IP_CLK) then
            if BUS2IP_RESET = '1' or IP2Shim_WrAck_int = '1' or IP2Shim_RdAck_int = '1' then
               shim2IP_CS   <= (others => '0');
               shim2IP_RdCE <= (others => '0');
               shim2IP_WrCE <= (others => '0');
               shim2IP_RNW  <= '0';
               Shim2IP_Addr <= (others => '0');
            else
               shim2IP_CS   <= shim2IP_CS_int  ;
               shim2IP_RdCE <= shim2IP_RdCE_int;
               shim2IP_WrCE <= shim2IP_WrCE_int;
               shim2IP_RNW  <= shim2IP_RNW_int;
               Shim2IP_Addr <= BUS2IP_Addr_reg;
            end if;
         end if;
      end process;


      ----------------------------------------------------------------------------
      -- Delay invalid response for rising edge detect
      ----------------------------------------------------------------------------
      DELAY_INVALID_RESPONSE : process (BUS2IP_CLK)
      begin

         if rising_edge(BUS2IP_CLK) then
            if BUS2IP_CS_reg = '1' then
               invalidAddrRspns_reg <= invalidAddrRspns;
            else
               invalidAddrRspns_reg <= '0';
            end if;
         end if;
      end process;



      ----------------------------------------------------------------------------
      -- Set invalid Request for Read transaction if it occured
      ----------------------------------------------------------------------------
      SET_INVALID_READ : process (BUS2IP_CLK)
      begin

         if rising_edge(BUS2IP_CLK) then
            if BUS2IP_RdCE_reg = '1' then
               --Pulse signal using rising edge detection
               invalidRdReq <= invalidAddrRspns and not invalidAddrRspns_reg;
            else
               invalidRdReq <= '0';
            end if;
         end if;
      end process;


      ----------------------------------------------------------------------------
      -- Set invalid Request for Write transaction if it occured
      ----------------------------------------------------------------------------
      SET_INVALID_WRITE : process (BUS2IP_CLK)
      begin

         if rising_edge(BUS2IP_CLK) then
            if BUS2IP_WrCE_reg = '1' then
               --Pulse signal using rising edge detection
               invalidWrReq <= invalidAddrRspns and not invalidAddrRspns_reg;
            else
               invalidWrReq <= '0';
            end if;
         end if;
      end process;

end rtl;



-------------------------------------------------------------------------------
-- tx_mem_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_mem_if.vhd
-- Version:         v1.00a
-- Description:     embedded ip transmit interface AXI Stream memory
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  tx_if.vhd
--                    tx_axistream_if.vhd
--          ->        tx_mem_if
--                    tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

--library lib_bmg_v1_0;
--use lib_bmg_v1_0.all;

Library xpm;
use xpm.vcomponents.all;

library work;
use work.tx_if_pack.all;




-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity tx_mem_if is
  generic (
    C_FAMILY               : string                      := "virtex6";

    -- Read Port - AXI Stream TxData
    c_TxD_write_width_a      : integer range   0 to 18     := 9;
    c_TxD_read_width_a       : integer range   0 to 18     := 9;
    c_TxD_write_depth_a      : integer range   0 to 32768  := 4096;
    c_TxD_read_depth_a       : integer range   0 to 32768  := 4096;
    c_TxD_addra_width        : integer range   0 to 15     := 10;
    c_TxD_wea_width          : integer range   0 to 2      := 2;
    -- Write Port - AXI Stream TxData
    c_TxD_write_width_b      : integer range  36 to 36     := 36;
    c_TxD_read_width_b       : integer range  36 to 36     := 36;
    c_TxD_write_depth_b      : integer range   0 to 8192   := 1024;
    c_TxD_read_depth_b       : integer range   0 to 8192   := 1024;
    c_TxD_addrb_width        : integer range   0 to 13     := 10;
    c_TxD_web_width          : integer range   0 to 4      := 4;

    -- Read Port - AXI Stream TxControl
    c_TxC_write_width_a      : integer range  36 to 36     := 36;
    c_TxC_read_width_a       : integer range  36 to 36     := 36;
    c_TxC_write_depth_a      : integer range   0 to 1024   := 1024;
    c_TxC_read_depth_a       : integer range   0 to 1024   := 1024;
    c_TxC_addra_width        : integer range   0 to 10     := 10;
    c_TxC_wea_width          : integer range   0 to 1      := 1;
    -- Write Port - AXI Stream TxControl
    c_TxC_write_width_b      : integer range   36 to 36    := 36;
    c_TxC_read_width_b       : integer range   36 to 36    := 36;
    c_TxC_write_depth_b      : integer range    0 to 1024  := 1024;
    c_TxC_read_depth_b       : integer range    0 to 1024  := 1024;
    c_TxC_addrb_width        : integer range    0 to 10    := 10;
    c_TxC_web_width          : integer range    0 to 1     := 1

  );
  port (
    -- Read Port - AXI Stream TxData
    TX_CLIENT_CLK             : in  std_logic;                                          --  Tx Client Clock
    reset2tx_client           : in  std_logic;                                          --  Reset
    Tx_Client_TxD_2_Mem_Din   : in  std_logic_vector(c_TxD_write_width_a-1 downto 0);   --  Tx Client Data Memory Wr Data
    Tx_Client_TxD_2_Mem_Addr  : in  std_logic_vector(c_TxD_addra_width-1   downto 0);   --  Tx Client Data Memory Address
    Tx_Client_TxD_2_Mem_En    : in  std_logic;                                          --  Tx Client Data Memory Enable
    Tx_Client_TxD_2_Mem_We    : in  std_logic_vector(c_TxD_wea_width-1     downto 0);   --  Tx Client Data Memory Wr Enable
    Tx_Client_TxD_2_Mem_Dout  : out std_logic_vector(c_TxD_read_width_a-1  downto 0);   --  Tx Client Data Memory Rd Data
    -- Write Port - AXI Stream TxData
    AXI_STR_TXD_ACLK          : in  std_logic;                                          --  AXI-Stream Tx Data Clock
    reset2axi_str_txd         : in  std_logic;                                          --  Reset
    Axi_Str_TxD_2_Mem_Din     : in  std_logic_vector(c_TxD_write_width_b-1 downto 0);   --  AXI-Stream Tx Data Memory Wr Data
    Axi_Str_TxD_2_Mem_Addr    : in  std_logic_vector(c_TxD_addrb_width-1   downto 0);   --  AXI-Stream Tx Data Memory Address
    Axi_Str_TxD_2_Mem_En      : in  std_logic;                                          --  AXI-Stream Tx Data Memory Enable
    Axi_Str_TxD_2_Mem_We      : in  std_logic_vector(c_TxD_web_width-1     downto 0);   --  AXI-Stream Tx Data Memory Wr Enable
    Axi_Str_TxD_2_Mem_Dout    : out std_logic_vector(c_TxD_read_width_b-1  downto 0);   --  AXI-Stream Tx Data Memory Rd Data

    -- Read Port - AXI Stream TxControl
    Tx_Client_TxC_2_Mem_Din   : in  std_logic_vector(c_TxC_write_width_a-1 downto 0);   --  Tx Client Control Memory Wr Data
    Tx_Client_TxC_2_Mem_Addr  : in  std_logic_vector(c_TxC_addra_width-1   downto 0);   --  Tx Client Control Memory Address
    Tx_Client_TxC_2_Mem_En    : in  std_logic;                                          --  Tx Client Control Memory Enable
    Tx_Client_TxC_2_Mem_We    : in  std_logic_vector(c_TxC_wea_width-1     downto 0);   --  Tx Client Control Memory Wr Enable
    Tx_Client_TxC_2_Mem_Dout  : out std_logic_vector(c_TxC_read_width_a-1  downto 0);   --  Tx Client Control Memory Rd Data
    -- Write Port - AXI Stream TxControl
    AXI_STR_TXC_ACLK          : in  std_logic;                                          --  AXI-Stream Tx Control Clock
    reset2axi_str_txc         : in  std_logic;                                          --  Reset
    Axi_Str_TxC_2_Mem_Din     : in  std_logic_vector(c_TxC_write_width_b-1 downto 0);   --  AXI-Stream Tx Control Memory Wr Data
    Axi_Str_TxC_2_Mem_Addr    : in  std_logic_vector(c_TxC_addrb_width-1   downto 0);   --  AXI-Stream Tx Control Memory Address
    Axi_Str_TxC_2_Mem_En      : in  std_logic;                                          --  AXI-Stream Tx Control Memory Enable
    Axi_Str_TxC_2_Mem_We      : in  std_logic_vector(c_TxC_web_width-1     downto 0);   --  AXI-Stream Tx Control Memory Wr Enable
    Axi_Str_TxC_2_Mem_Dout    : out std_logic_vector(c_TxC_read_width_b-1  downto 0)    --  AXI-Stream Tx Control Memory Rd Data
  );

end tx_mem_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture imp of tx_mem_if is

begin

-- XPM Memory between AXI Stream Interface and Tx Client Interface

-- Start of xpm_memory_tdpram_inst instance declaration

TXD_MEM : xpm_memory_tdpram
  generic map (

    -- Common module generics
    MEMORY_SIZE             => c_TxD_write_width_a*c_TxD_write_depth_a,            --positive integer
    MEMORY_PRIMITIVE        => "block",          --string; "auto", "distributed", "block" or "ultra" ;
    CLOCKING_MODE           => "independent_clock",  --string; "common_clock", "independent_clock" 
    MEMORY_INIT_FILE        => "none",          --string; "none" or "<filename>.mem" 
    MEMORY_INIT_PARAM       => "",              --string;
    USE_MEM_INIT            => 1,               --integer; 0,1
    WAKEUP_TIME             => "disable_sleep", --string; "disable_sleep" or "use_sleep_pin" 
    MESSAGE_CONTROL         => 0,               --integer;
    ECC_MODE                => "no_ecc",        --string; "no_ecc", "encode_only", "decode_only" or "both_encode_and_decode" 
    AUTO_SLEEP_TIME         => 0,               --Do not Change
    USE_EMBEDDED_CONSTRAINT => 0,               --integer: 0,1
    MEMORY_OPTIMIZATION     => "true",          --string; "true", "false" 

    -- Port A module generics
    WRITE_DATA_WIDTH_A      => c_TxD_write_width_a,              --positive integer
    READ_DATA_WIDTH_A       => c_TxD_read_width_a,              --positive integer
    BYTE_WRITE_WIDTH_A      => c_TxD_write_width_a/c_TxD_wea_width,              --integer; 8, 9, or WRITE_DATA_WIDTH_A value
    ADDR_WIDTH_A            => c_TxD_addra_width,               --positive integer
    READ_RESET_VALUE_A      => "0",             --string
    READ_LATENCY_A          => 1,               --non-negative integer
    WRITE_MODE_A            => "write_first",     --string; "write_first", "read_first", "no_change" 

    -- Port B module generics
    WRITE_DATA_WIDTH_B      => c_TxD_write_width_b,              --positive integer
    READ_DATA_WIDTH_B       => c_TxD_read_width_b,              --positive integer
    BYTE_WRITE_WIDTH_B      => c_TxD_write_width_b/c_TxD_web_width,              --integer; 8, 9, or WRITE_DATA_WIDTH_B value
    ADDR_WIDTH_B            => c_TxD_addrb_width,               --positive integer
    READ_RESET_VALUE_B      => "0",             --string
    READ_LATENCY_B          => 1,               --non-negative integer
    WRITE_MODE_B            => "write_first"      --string; "write_first", "read_first", "no_change" 
  )
  port map (

    -- Common module ports
    sleep                   => '0',

    -- Port A module ports
    clka                    => TX_CLIENT_CLK,
    rsta                    => reset2tx_client,
    ena                     => Tx_Client_TxD_2_Mem_En,
    regcea                  => '0',
    wea                     => Tx_Client_TxD_2_Mem_We, 
    addra                   => Tx_Client_TxD_2_Mem_Addr,
    dina                    => Tx_Client_TxD_2_Mem_Din,
    injectsbiterra          => '0',
    injectdbiterra          => '0',
    douta                   => Tx_Client_TxD_2_Mem_Dout,
    sbiterra                => open,
    dbiterra                => open,

    -- Port B module ports
    clkb                    => AXI_STR_TXD_ACLK,
    rstb                    => reset2axi_str_txd,
    enb                     => Axi_Str_TxD_2_Mem_En,
    regceb                  => '0',
    web                     => Axi_Str_TxD_2_Mem_We, 
    addrb                   => Axi_Str_TxD_2_Mem_Addr,
    dinb                    => Axi_Str_TxD_2_Mem_Din,
    injectsbiterrb          => '0',
    injectdbiterrb          => '0',
    doutb                   => Axi_Str_TxD_2_Mem_Dout,
    sbiterrb                => open,
    dbiterrb                => open
  );

-- End of xpm_memory_tdpram_inst instance declaration

--  TXD_MEM : entity lib_bmg_v1_0.blk_mem_gen_wrapper(implementation)
--  --BRAM between AXI Stream Interface and Tx Client Interface
--  generic map(
--    c_family                 => C_FAMILY,
--    c_xdevicefamily          => C_FAMILY,
--
--    -- Selection between BMG and XPM
--    bmg_xpm_sel              => 1,
--    -- Memory Specific Configurations
--    c_mem_type               => 2,
--       -- This wrapper only supports the True Dual Port RAM
--       -- 0: Single Port RAM
--       -- 1: Simple Dual Port RAM
--       -- 2: True Dual Port RAM
--       -- 3: Single Port Rom
--       -- 4: Dual Port RAM
--    c_algorithm              => 1,
--       -- 0: Selectable Primative
--       -- 1: Minimum Area
--    c_prim_type              => 3,
--       -- 0: ( 1-bit wide)
--       -- 1: ( 2-bit wide)
--       -- 2: ( 4-bit wide)
--       -- 3: ( 9-bit wide)
--       -- 4: (18-bit wide)
--       -- 5: (36-bit wide)
--       -- 6: (72-bit wide, single port only)
--    c_byte_size              => 9,   -- 8 or 9
--
--    -- Simulation Behavior Options
--    c_sim_collision_check    => "NONE",
--       -- "None"
--       -- "Generate_X"
--       -- "All"
--       -- "Warnings_only"
--    c_common_clk             => 0,   -- 0, 1
--    c_disable_warn_bhv_coll  => 0,   -- 0, 1
--    c_disable_warn_bhv_range => 0,   -- 0, 1
--
--    -- Initialization Configuration Options
--    c_load_init_file         => 0,
--    c_init_file_name         => "none",
--    c_use_default_data       => 0,   -- 0, 1
--    c_default_data           => "0", -- "..."
--
--    -- Port A Specific Configurations - 8bit bus
--    c_has_mem_output_regs_a  => 0,   -- 0, 1
--    c_has_mux_output_regs_a  => 0,   -- 0, 1
--    c_write_width_a          => c_TxD_write_width_a,  -- 1 to 1152
--    c_read_width_a           => c_TxD_read_width_a,  -- 1 to 1152
--    c_write_depth_a          => c_TxD_write_depth_a,  -- 2 to 9011200
--    c_read_depth_a           => c_TxD_read_depth_a,  -- 2 to 9011200
--    c_addra_width            => c_TxD_addra_width,   -- 1 to 24
--    c_write_mode_a           => "WRITE_FIRST",  -- Need to use "WRITE_FIRST" instead of "NO CHANGE" to use byte write enable
--       -- "Write_First"
--       -- "Read_first"
--       -- "No_Change"
--    c_has_ena                => 1,   -- 0, 1
--    c_has_regcea             => 0,   -- 0, 1
--    c_has_ssra               => 1,   -- 0, 1
--    c_sinita_val             => "0", --"..."
--    c_use_byte_wea           => 1,   -- 0, 1
--    c_wea_width              => c_TxD_wea_width,   -- 1 to 128
--
--    -- Port B Specific Configurations - 32bit bus
--    c_has_mem_output_regs_b  => 0,   -- 0, 1
--    c_has_mux_output_regs_b  => 0,   -- 0, 1
--    c_write_width_b          => c_TxD_write_width_b,  -- 1 to 1152
--    c_read_width_b           => c_TxD_read_width_b,  -- 1 to 1152
--    c_write_depth_b          => c_TxD_write_depth_b,  -- 2 to 9011200
--    c_read_depth_b           => c_TxD_read_depth_b,   -- 2 to 9011200
--    c_addrb_width            => c_TxD_addrb_width,   -- 1 to 24
--    c_write_mode_b           => "WRITE_FIRST",  -- Need to use "WRITE_FIRST" instead of "NO CHANGE" to use byte write enable
--       -- "Write_First"
--       -- "Read_first"
--       -- "No_Change"
--    c_has_enb                => 1,   -- 0, 1
--    c_has_regceb             => 0,   -- 0, 1
--    c_has_ssrb               => 1,   -- 0, 1
--    c_sinitb_val             => "0", -- "..."
--    c_use_byte_web           => 1,   -- 0, 1
--    c_web_width              => c_TxD_web_width,   -- 1 to 128
--
--    -- Other Miscellaneous Configurations
--    c_mux_pipeline_stages    => 0,   -- 0, 1, 2, 3
--       -- The number of pipeline stages within the MUX
--       --    for both Port A and Port B
--    c_use_ecc                => 0,
--       -- See DS512 for the limited core option selections for ECC support
--    c_use_ramb16bwer_rst_bhv => 0    --0, 1
--  )
--  port map  (
--    -- Read Port
--    clka    => TX_CLIENT_CLK,            --: in  std_logic;
--    ssra    => reset2tx_client,          --: in  std_logic := '0';
--    dina    => Tx_Client_TxD_2_Mem_Din,  --: in  std_logic_vector(c_write_width_a-1 downto 0) := (OTHERS => '0');
--    addra   => Tx_Client_TxD_2_Mem_Addr, --: in  std_logic_vector(c_addra_width-1   downto 0);
--    ena     => Tx_Client_TxD_2_Mem_En,   --: in  std_logic := '1';
--    regcea  => '0',                      --: in  std_logic := '1';
--    wea     => Tx_Client_TxD_2_Mem_We,   --: in  std_logic_vector(c_wea_width-1     downto 0) := (OTHERS => '0');
--    douta   => Tx_Client_TxD_2_Mem_Dout, --: out std_logic_vector(c_read_width_a-1  downto 0);
--    --  Write Port
--    clkb    => AXI_STR_TXD_ACLK,         --: in  std_logic := '0';
--    ssrb    => reset2axi_str_txd,        --: in  std_logic := '0';
--    dinb    => Axi_Str_TxD_2_Mem_Din,    --: in  std_logic_vector(c_write_width_b-1 downto 0) := (OTHERS => '0');
--    addrb   => Axi_Str_TxD_2_Mem_Addr,   --: in  std_logic_vector(c_addrb_width-1   downto 0) := (OTHERS => '0');
--    enb     => Axi_Str_TxD_2_Mem_En,     --: in  std_logic := '1';
--    regceb  => '0',                      --: in  std_logic := '1';
--    web     => Axi_Str_TxD_2_Mem_We,     --: in  std_logic_vector(c_web_width-1     downto 0) := (OTHERS => '0');
--    doutb   => Axi_Str_TxD_2_Mem_Dout,                 --: out std_logic_vector(c_read_width_b-1  downto 0);
--
--    dbiterr => open,                 --: out std_logic;
--                                     -- Double bit error that that cannot be auto corrected by ECC
--    sbiterr => open                  --: out std_logic
--
--  );

-- XPM Memory between AXI Stream Interface and Tx Client Interface

-- Start of xpm_memory_tdpram_inst instance declaration

TXC_MEM: xpm_memory_tdpram
  generic map (

    -- Common module generics
    MEMORY_SIZE             => c_TxC_write_width_a*c_TxC_write_depth_a,            --positive integer
    MEMORY_PRIMITIVE        => "block",          --string; "auto", "distributed", "block" or "ultra" ;
    CLOCKING_MODE           => "independent_clock",  --string; "common_clock", "independent_clock" 
    MEMORY_INIT_FILE        => "none",          --string; "none" or "<filename>.mem" 
    MEMORY_INIT_PARAM       => "",              --string;
    USE_MEM_INIT            => 1,               --integer; 0,1
    WAKEUP_TIME             => "disable_sleep", --string; "disable_sleep" or "use_sleep_pin" 
    MESSAGE_CONTROL         => 0,               --integer;
    ECC_MODE                => "no_ecc",        --string; "no_ecc", "encode_only", "decode_only" or "both_encode_and_decode" 
    AUTO_SLEEP_TIME         => 0,               --Do not Change
    USE_EMBEDDED_CONSTRAINT => 0,               --integer: 0,1
    MEMORY_OPTIMIZATION     => "true",          --string; "true", "false" 

    -- Port A module generics
    WRITE_DATA_WIDTH_A      => c_TxC_write_width_a,              --positive integer
    READ_DATA_WIDTH_A       => c_TxC_read_width_a,              --positive integer
    BYTE_WRITE_WIDTH_A      => c_TxC_write_width_a/c_TxC_wea_width,              --integer; 8, 9, or WRITE_DATA_WIDTH_A value
    ADDR_WIDTH_A            => c_TxC_addra_width,               --positive integer
    READ_RESET_VALUE_A      => "0",             --string
    READ_LATENCY_A          => 1,               --non-negative integer
    WRITE_MODE_A            => "no_change",     --string; "write_first", "read_first", "no_change" 

    -- Port B module generics
    WRITE_DATA_WIDTH_B      => c_TxC_write_width_b,              --positive integer
    READ_DATA_WIDTH_B       => c_TxC_read_width_b,              --positive integer
    BYTE_WRITE_WIDTH_B      => c_TxC_write_width_b/c_TxC_web_width,              --integer; 8, 9, or WRITE_DATA_WIDTH_B value
    ADDR_WIDTH_B            => c_TxC_addrb_width,               --positive integer
    READ_RESET_VALUE_B      => "0",             --string
    READ_LATENCY_B          => 1,               --non-negative integer
    WRITE_MODE_B            => "no_change"      --string; "write_first", "read_first", "no_change" 
  )
  port map (

    -- Common module ports
    sleep                   => '0',

    -- Port A module ports
    clka                    => TX_CLIENT_CLK,
    rsta                    => reset2tx_client,
    ena                     => Tx_Client_TxC_2_Mem_En,
    regcea                  => '0',
    wea                     => Tx_Client_TxC_2_Mem_We,
    addra                   => Tx_Client_TxC_2_Mem_Addr,
    dina                    => Tx_Client_TxC_2_Mem_Din,
    injectsbiterra          => '0',
    injectdbiterra          => '0',
    douta                   => Tx_Client_TxC_2_Mem_Dout,
    sbiterra                => open,
    dbiterra                => open,

    -- Port B module ports
    clkb                    => AXI_STR_TXC_ACLK,
    rstb                    => reset2axi_str_txc,
    enb                     => Axi_Str_TxC_2_Mem_En,
    regceb                  => '0',
    web                     => Axi_Str_TxC_2_Mem_We,
    addrb                   => Axi_Str_TxC_2_Mem_Addr,
    dinb                    => Axi_Str_TxC_2_Mem_Din,
    injectsbiterrb          => '0',
    injectdbiterrb          => '0',
    doutb                   => Axi_Str_TxC_2_Mem_Dout,
    sbiterrb                => open,
    dbiterrb                => open
  );

-- End of xpm_memory_tdpram_inst instance declaration

--  TXC_MEM : entity lib_bmg_v1_0.blk_mem_gen_wrapper(implementation)
--  --BRAM between AXI Stream Interface and Tx Client Interface
--  generic map(
--    c_family                 => C_FAMILY,
--    c_xdevicefamily          => C_FAMILY,
--
--    -- Selection between BMG and XPM
--    bmg_xpm_sel              => 0,
--    -- Memory Specific Configurations
--    c_mem_type               => 2,
--       -- This wrapper only supports the True Dual Port RAM
--       -- 0: Single Port RAM
--       -- 1: Simple Dual Port RAM
--       -- 2: True Dual Port RAM
--       -- 3: Single Port Rom
--       -- 4: Dual Port RAM
--    c_algorithm              => 1,
--       -- 0: Selectable Primative
--       -- 1: Minimum Area
--    c_prim_type              => 3,
--       -- 0: ( 1-bit wide)
--       -- 1: ( 2-bit wide)
--       -- 2: ( 4-bit wide)
--       -- 3: ( 9-bit wide)
--       -- 4: (18-bit wide)
--       -- 5: (36-bit wide)
--       -- 6: (72-bit wide, single port only)
--    c_byte_size              => 9,   -- 8 or 9
--
--    -- Simulation Behavior Options
--    c_sim_collision_check    => "NONE",
--       -- "None"
--       -- "Generate_X"
--       -- "All"
--       -- "Warnings_only"
--    c_common_clk             => 0,   -- 0, 1
--    c_disable_warn_bhv_coll  => 0,   -- 0, 1
--    c_disable_warn_bhv_range => 0,   -- 0, 1
--
--    -- Initialization Configuration Options
--    c_load_init_file         => 0,
--    c_init_file_name         => "none",
--    c_use_default_data       => 1,   -- 0, 1
--    c_default_data           => "0", -- "..."
--
--    -- Port A Specific Configurations - 8bit bus
--    c_has_mem_output_regs_a  => 0,   -- 0, 1
--    c_has_mux_output_regs_a  => 0,   -- 0, 1
--    c_write_width_a          => c_TxC_write_width_a,  -- 1 to 1152
--    c_read_width_a           => c_TxC_read_width_a,  -- 1 to 1152
--    c_write_depth_a          => c_TxC_write_depth_a,  -- 2 to 9011200
--    c_read_depth_a           => c_TxC_read_depth_a,  -- 2 to 9011200
--    c_addra_width            => c_TxC_addra_width,   -- 1 to 24
--    c_write_mode_a           => "NO_CHANGE",
--       -- "Write_First"
--       -- "Read_first"
--       -- "No_Change"
--    c_has_ena                => 1,   -- 0, 1
--    c_has_regcea             => 0,   -- 0, 1
--    c_has_ssra               => 1,   -- 0, 1
--    c_sinita_val             => "0", --"..."
--    c_use_byte_wea           => 0,   -- 0, 1
--    c_wea_width              => c_TxC_wea_width,   -- 1 to 128
--
--    -- Port B Specific Configurations - 32bit bus
--    c_has_mem_output_regs_b  => 0,   -- 0, 1
--    c_has_mux_output_regs_b  => 0,   -- 0, 1
--    c_write_width_b          => c_TxC_write_width_b,  -- 1 to 1152
--    c_read_width_b           => c_TxC_read_width_b,  -- 1 to 1152
--    c_write_depth_b          => c_TxC_write_depth_b,  -- 2 to 9011200
--    c_read_depth_b           => c_TxC_read_depth_b,   -- 2 to 9011200
--    c_addrb_width            => c_TxC_addrb_width,   -- 1 to 24
--    c_write_mode_b           => "NO_CHANGE",
--       -- "Write_First"
--       -- "Read_first"
--       -- "No_Change"
--    c_has_enb                => 1,   -- 0, 1
--    c_has_regceb             => 0,   -- 0, 1
--    c_has_ssrb               => 1,   -- 0, 1
--    c_sinitb_val             => "0", -- "..."
--    c_use_byte_web           => 0,   -- 0, 1
--    c_web_width              => c_TxC_web_width,   -- 1 to 128
--
--    -- Other Miscellaneous Configurations
--    c_mux_pipeline_stages    => 0,   -- 0, 1, 2, 3
--       -- The number of pipeline stages within the MUX
--       --    for both Port A and Port B
--    c_use_ecc                => 0,
--       -- See DS512 for the limited core option selections for ECC support
--    c_use_ramb16bwer_rst_bhv => 0    --0, 1
--  )
--  port map  (
--    -- Read Port
--    clka    => TX_CLIENT_CLK,            --: in  std_logic;
--    ssra    => reset2tx_client,          --: in  std_logic := '0';
--    dina    => Tx_Client_TxC_2_Mem_Din,  --: in  std_logic_vector(c_write_width_a-1 downto 0) := (OTHERS => '0');
--    addra   => Tx_Client_TxC_2_Mem_Addr, --: in  std_logic_vector(c_addra_width-1   downto 0);
--    ena     => Tx_Client_TxC_2_Mem_En,   --: in  std_logic := '1';
--    regcea  => '0',                      --: in  std_logic := '1';
--    wea     => Tx_Client_TxC_2_Mem_We,   --: in  std_logic_vector(c_wea_width-1     downto 0) := (OTHERS => '0');
--    douta   => Tx_Client_TxC_2_Mem_Dout, --: out std_logic_vector(c_read_width_a-1  downto 0);
--    --  Write Port
--    clkb    => AXI_STR_TXC_ACLK,         --: in  std_logic := '0';
--    ssrb    => reset2axi_str_txc,        --: in  std_logic := '0';
--    dinb    => Axi_Str_TxC_2_Mem_Din,    --: in  std_logic_vector(c_write_width_b-1 downto 0) := (OTHERS => '0');
--    addrb   => Axi_Str_TxC_2_Mem_Addr,   --: in  std_logic_vector(c_addrb_width-1   downto 0) := (OTHERS => '0');
--    enb     => Axi_Str_TxC_2_Mem_En,     --: in  std_logic := '1';
--    regceb  => '0',                      --: in  std_logic := '1';
--    web     => Axi_Str_TxC_2_Mem_We,     --: in  std_logic_vector(c_web_width-1     downto 0) := (OTHERS => '0');
--    doutb   => Axi_Str_TxC_2_Mem_Dout,   --: out std_logic_vector(c_read_width_b-1  downto 0);
--
--    dbiterr => open,                 --: out std_logic;
--                                     -- Double bit error that that cannot be auto corrected by ECC
--    sbiterr => open                  --: out std_logic
--
--  );

end imp;


------------------------------------------------------------------------------
-- rx_mem_if.vhd
------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        rx_mem_if.vhd
-- Version:         v1.00a
-- Description:     Receive interface between AXIStream and Temac
--
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--                  rx_if.vhd
--                    rx_axistream_if.vhd
--          ->        rx_mem_if
--                    rx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MSH
--
--  MSH     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Libraries used;
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

--library lib_bmg_v1_0;
--use lib_bmg_v1_0.all;

Library xpm;
use xpm.vcomponents.all;

library work;
use work.rx_if_pack.all;

-------------------------------------------------------------------------------
-- Definition of Generics :
-------------------------------------------------------------------------------
--
--  C_FAMILY              -- Xilinx FPGA Family
--  C_RXD_MEM_ADDR_WIDTH           --
--  C_RXD_MEM_BYTES
--  C_RXS_MEM_ADDR_WIDTH           --
--  C_RXS_MEM_BYTES
--
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Definition of Ports :
-------------------------------------------------------------------------------
--
--  AXI_STR_RXD_ACLK
--  AXI_STR_RXD_DPMEM_WR_DATA
--  AXI_STR_RXD_DPMEM_RD_DATA
--  AXI_STR_RXD_DPMEM_WR_EN
--  AXI_STR_RXD_DPMEM_ADDR
--
--  AXI_STR_RXS_ACLK
--  AXI_STR_RXS_DPMEM_WR_DATA
--  AXI_STR_RXS_DPMEM_RD_DATA
--  AXI_STR_RXS_DPMEM_WR_EN
--  AXI_STR_RXS_DPMEM_ADDR
--
--  RX_CLIENT_CLK
--  RX_CLIENT_CLK_ENBL
--  RX_CLIENT_RXD_DPMEM_WR_DATA
--  RX_CLIENT_RXD_DPMEM_RD_DATA
--  RX_CLIENT_RXD_DPMEM_WR_EN
--  RX_CLIENT_RXD_DPMEM_ADDR
--  RESET2RX_CLIENT
--
--  RX_CLIENT_RXS_DPMEM_WR_DATA
--  RX_CLIENT_RXS_DPMEM_RD_DATA
--  RX_CLIENT_RXS_DPMEM_WR_EN
--  RX_CLIENT_RXS_DPMEM_ADDR
--
-------------------------------------------------------------------------------
----                  Entity Section
-------------------------------------------------------------------------------

entity rx_mem_if is
  generic (
    C_RXD_MEM_BYTES      : integer    := 4096;
    C_RXD_MEM_ADDR_WIDTH : integer    := 10;
    C_RXS_MEM_BYTES      : integer    := 4096;
    C_RXS_MEM_ADDR_WIDTH : integer    := 10;
    C_FAMILY             : string     := "virtex6"
  );

  port    (
    AXI_STR_RXD_ACLK            : in  std_logic;                                        --  AXI-Stream Receive Data Clock
    AXI_STR_RXD_DPMEM_WR_DATA   : in  std_logic_vector(35 downto 0);                    --  AXI-Stream Receive Data Write Data
    AXI_STR_RXD_DPMEM_RD_DATA   : out std_logic_vector(35 downto 0);                    --  AXI-Stream Receive Data Read Data
    AXI_STR_RXD_DPMEM_WR_EN     : in  std_logic_vector(0 downto 0);                     --  AXI-Stream Receive Data Write Enable
    AXI_STR_RXD_DPMEM_ADDR      : in  std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  AXI-Stream Receive Data Address
    RESET2AXI_STR_RXD           : in  std_logic;                                        --  AXI-Stream Receive Data Rese

    AXI_STR_RXS_ACLK            : in  std_logic;                                        --  AXI-Stream Receive Status Clock
    AXI_STR_RXS_DPMEM_WR_DATA   : in  std_logic_vector(35 downto 0);                    --  AXI-Stream Receive Status Write Data
    AXI_STR_RXS_DPMEM_RD_DATA   : out std_logic_vector(35 downto 0);                    --  AXI-Stream Receive Status Read Data
    AXI_STR_RXS_DPMEM_WR_EN     : in  std_logic_vector(0 downto 0);                     --  AXI-Stream Receive Status Write Enable
    AXI_STR_RXS_DPMEM_ADDR      : in  std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  AXI-Stream Receive Status Address
    RESET2AXI_STR_RXS           : in  std_logic;                                        --  AXI-Stream Receive Status Rese

    RX_CLIENT_CLK               : in  std_logic;                                        --  Receive MAC Clock
    RX_CLIENT_CLK_ENBL          : in  std_logic;                                        --  Receive MAC Clock Enable
    RX_CLIENT_RXD_DPMEM_WR_DATA : in  std_logic_vector(35 downto 0);                    --  Receive MAC Data Memory Write Data
    RX_CLIENT_RXD_DPMEM_RD_DATA : out std_logic_vector(35 downto 0);                    --  Receive MAC Data Memory Read Data
    RX_CLIENT_RXD_DPMEM_WR_EN   : in  std_logic_vector(0 downto 0);                     --  Receive MAC Data Memory Write Enable
    RX_CLIENT_RXD_DPMEM_ADDR    : in  std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);  --  Receive MAC Data Memory Address

    RX_CLIENT_RXS_DPMEM_WR_DATA : in  std_logic_vector(35 downto 0);                    --  Receive MAC Status Memory Write Data
    RX_CLIENT_RXS_DPMEM_RD_DATA : out std_logic_vector(35 downto 0);                    --  Receive MAC Status Memory Read Data
    RX_CLIENT_RXS_DPMEM_WR_EN   : in  std_logic_vector(0 downto 0);                     --  Receive MAC Status Memory Write Enable
    RX_CLIENT_RXS_DPMEM_ADDR    : in  std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);  --  Receive MAC Status Memory Address
    RESET2RX_CLIENT         : in  std_logic                                             --  Receive MAC Reset
  );
end rx_mem_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of rx_mem_if is

function log2(x : natural) return integer is
  variable i  : integer := 0;
  variable val: integer := 1;
begin
  if x = 0 then return 0;
  else
    for j in 0 to 29 loop -- for loop for XST 
      if val >= x then null;
      else
        i := i+1;
        val := val*2;
      end if;
    end loop;
  -- synthesis translate_off
    assert val >= x
      report "Function log2 received argument larger" &
             " than its capability of 2^30. "
      severity failure;
  -- synthesis translate_on
    return i;
  end if;
end function log2;

------------------------------------------------------------------------------
-- Constant Declarations
------------------------------------------------------------------------------


------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------
signal rx_client_rxs_dpmem_wr_data_d1 :  std_logic_vector(35 downto 0);
signal rx_client_rxs_dpmem_wr_en_d1   :  std_logic_vector(0 downto 0);
signal rx_client_rxs_dpmem_addr_d1    :  std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal rx_client_rxd_dpmem_wr_data_d1 :  std_logic_vector(35 downto 0);
signal rx_client_rxd_dpmem_wr_en_d1   :  std_logic_vector(0 downto 0);
signal rx_client_rxd_dpmem_addr_d1    :  std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);

signal rx_client_clk_enbl_d1          :  std_logic;


begin

  PIPELINE_RXSMEMREG : process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        rx_client_rxs_dpmem_wr_data_d1 <= (others => '0');
        rx_client_rxs_dpmem_wr_en_d1   <= (others => '0');
        rx_client_rxs_dpmem_addr_d1    <= (others => '0');
        rx_client_clk_enbl_d1          <= '0';
      else
        rx_client_rxs_dpmem_wr_data_d1 <= RX_CLIENT_RXS_DPMEM_WR_DATA;
        rx_client_rxs_dpmem_wr_en_d1   <= RX_CLIENT_RXS_DPMEM_WR_EN;
        rx_client_rxs_dpmem_addr_d1    <= RX_CLIENT_RXS_DPMEM_ADDR;
        rx_client_clk_enbl_d1          <= RX_CLIENT_CLK_ENBL;
      end if;
    end if;
  end process;

  PIPELINE_RXDMEMREG : process (RX_CLIENT_CLK)
  begin
    if rising_edge(RX_CLIENT_CLK) then
      if RESET2RX_CLIENT = '1' then
        rx_client_rxd_dpmem_wr_data_d1 <= (others => '0');
        rx_client_rxd_dpmem_wr_en_d1 <= (others => '0');
        rx_client_rxd_dpmem_addr_d1 <= (others => '0');
      else
        rx_client_rxd_dpmem_wr_data_d1 <= RX_CLIENT_RXD_DPMEM_WR_DATA;
        rx_client_rxd_dpmem_wr_en_d1 <= RX_CLIENT_RXD_DPMEM_WR_EN;
        rx_client_rxd_dpmem_addr_d1 <= RX_CLIENT_RXD_DPMEM_ADDR;
      end if;
    end if;
  end process;

-- Start of xpm_memory_tdpram_inst instance declaration

I_RXD_MEM: xpm_memory_tdpram
  generic map (

    -- Common module generics
    MEMORY_SIZE             => 36*(C_RXD_MEM_BYTES/4),            --positive integer
    MEMORY_PRIMITIVE        => "block",          --string; "auto", "distributed", "block" or "ultra" ;
    CLOCKING_MODE           => "independent_clock",  --string; "common_clock", "independent_clock" 
    MEMORY_INIT_FILE        => "none",          --string; "none" or "<filename>.mem" 
    MEMORY_INIT_PARAM       => "",              --string;
    USE_MEM_INIT            => 1,               --integer; 0,1
    WAKEUP_TIME             => "disable_sleep", --string; "disable_sleep" or "use_sleep_pin" 
    MESSAGE_CONTROL         => 0,               --integer;
    ECC_MODE                => "no_ecc",        --string; "no_ecc", "encode_only", "decode_only" or "both_encode_and_decode" 
    AUTO_SLEEP_TIME         => 0,               --Do not Change
    USE_EMBEDDED_CONSTRAINT => 0,               --integer: 0,1
    MEMORY_OPTIMIZATION     => "true",          --string; "true", "false" 

    -- Port A module generics
    WRITE_DATA_WIDTH_A      => 36,              --positive integer
    READ_DATA_WIDTH_A       => 36,              --positive integer
    BYTE_WRITE_WIDTH_A      => 36,              --integer; 8, 9, or WRITE_DATA_WIDTH_A value
    ADDR_WIDTH_A            => (log2(C_RXD_MEM_BYTES/4)),               --positive integer
    READ_RESET_VALUE_A      => "0",             --string
    READ_LATENCY_A          => 1,               --non-negative integer
    WRITE_MODE_A            => "no_change",     --string; "write_first", "read_first", "no_change" 

    -- Port B module generics
    WRITE_DATA_WIDTH_B      => 36,              --positive integer
    READ_DATA_WIDTH_B       => 36,              --positive integer
    BYTE_WRITE_WIDTH_B      => 36,              --integer; 8, 9, or WRITE_DATA_WIDTH_B value
    ADDR_WIDTH_B            => (log2(C_RXD_MEM_BYTES/4)),               --positive integer
    READ_RESET_VALUE_B      => "0",             --string
    READ_LATENCY_B          => 1,               --non-negative integer
    WRITE_MODE_B            => "no_change"      --string; "write_first", "read_first", "no_change" 
  )
  port map (

    -- Common module ports
    sleep                   => '0',

    -- Port A module ports
    clka                    => RX_CLIENT_CLK,
    rsta                    => RESET2RX_CLIENT,
    ena                     => rx_client_clk_enbl_d1,
    regcea                  => '0',
    wea                     => rx_client_rxd_dpmem_wr_en_d1,
    addra                   => rx_client_rxd_dpmem_addr_d1,
    dina                    => rx_client_rxd_dpmem_wr_data_d1,
    injectsbiterra          => '0',
    injectdbiterra          => '0',
    douta                   => RX_CLIENT_RXD_DPMEM_RD_DATA,
    sbiterra                => open,
    dbiterra                => open,

    -- Port B module ports
    clkb                    => AXI_STR_RXD_ACLK,
    rstb                    => RESET2AXI_STR_RXD,
    enb                     => '1',
    regceb                  => '0',
    web                     => AXI_STR_RXD_DPMEM_WR_EN,
    addrb                   => AXI_STR_RXD_DPMEM_ADDR,
    dinb                    => AXI_STR_RXD_DPMEM_WR_DATA,
    injectsbiterrb          => '0',
    injectdbiterrb          => '0',
    doutb                   => AXI_STR_RXD_DPMEM_RD_DATA,
    sbiterrb                => open,
    dbiterrb                => open
  );

-- End of xpm_memory_tdpram_inst instance declaration
-- I_RXD_MEM : entity lib_bmg_v1_0.blk_mem_gen_wrapper
--   generic map(
--      c_family                 => C_FAMILY,
--      c_xdevicefamily          => C_FAMILY,
--      -- Selection between BMG and XPM
--      bmg_xpm_sel              => 0,
--      -- Memory Specific Configurations
--      c_mem_type               => 2,
--         -- This wrapper only supports the True Dual Port RAM
--         -- 0: Single Port RAM
--         -- 1: Simple Dual Port RAM
--         -- 2: True Dual Port RAM
--         -- 3: Single Port Rom
--         -- 4: Dual Port RAM
--      c_algorithm              => 1,
--         -- 0: Selectable Primative
--         -- 1: Minimum Area
--      c_prim_type              => 1,
--         -- 0: ( 1-bit wide)
--         -- 1: ( 2-bit wide)
--         -- 2: ( 4-bit wide)
--         -- 3: ( 9-bit wide)
--         -- 4: (18-bit wide)
--         -- 5: (36-bit wide)
--         -- 6: (72-bit wide, single port only)
--      c_byte_size              => 9,   -- 8 or 9
--
--      -- Simulation Behavior Options
--      c_sim_collision_check    => "NONE",
--         -- "None"
--         -- "Generate_X"
--         -- "All"
--         -- "Warnings_only"
--      c_common_clk             => 0,   -- 0, 1
--      c_disable_warn_bhv_coll  => 0,   -- 0, 1
--      c_disable_warn_bhv_range => 0,   -- 0, 1
--
--      -- Initialization Configuration Options
--      c_load_init_file         => 0,
--      c_init_file_name         => "none",
--      c_use_default_data       => 0,   -- 0, 1
--      c_default_data           => "0", -- "..."
--
--      -- Port A Specific Configurations
--      c_has_mem_output_regs_a  => 0,   -- 0, 1
--      c_has_mux_output_regs_a  => 0,   -- 0, 1
--      c_write_width_a          => 36,  -- 1 to 1152
--      c_read_width_a           => 36,  -- 1 to 1152
--      c_write_depth_a          => (C_RXD_MEM_BYTES/4),  -- 2 to 9011200
--      c_read_depth_a           => (C_RXD_MEM_BYTES/4),  -- 2 to 9011200
--      c_addra_width            => (log2(C_RXD_MEM_BYTES/4)),   -- 1 to 24
--      c_write_mode_a           => "NO_CHANGE",
--         -- "Write_First"
--         -- "Read_first"
--         -- "No_Change"
--      c_has_ena                => 1,   -- 0, 1
--      c_has_regcea             => 0,   -- 0, 1
--      c_has_ssra               => 0,   -- 0, 1
--      c_sinita_val             => "0", --"..."
--      c_use_byte_wea           => 0,   -- 0, 1
--      c_wea_width              => 1,   -- 1 to 128
--
--      -- Port B Specific Configurations
--      c_has_mem_output_regs_b  => 0,   -- 0, 1
--      c_has_mux_output_regs_b  => 0,   -- 0, 1
--      c_write_width_b          => 36,  -- 1 to 1152
--      c_read_width_b           => 36,  -- 1 to 1152
--      c_write_depth_b          => (C_RXD_MEM_BYTES/4),  -- 2 to 9011200
--      c_read_depth_b           => (C_RXD_MEM_BYTES/4),   -- 2 to 9011200
--      c_addrb_width            => (log2(C_RXD_MEM_BYTES/4)),   -- 1 to 24
--      c_write_mode_b           => "NO_CHANGE",
--         -- "Write_First"
--         -- "Read_first"
--         -- "No_Change"
--      c_has_enb                => 0,   -- 0, 1
--      c_has_regceb             => 0,   -- 0, 1
--      c_has_ssrb               => 0,   -- 0, 1
--      c_sinitb_val             => "0", -- "..."
--      c_use_byte_web           => 0,   -- 0, 1
--      c_web_width              => 1,   -- 1 to 128
--
--      -- Other Miscellaneous Configurations
--      c_mux_pipeline_stages    => 0,   -- 0, 1, 2, 3
--         -- The number of pipeline stages within the MUX
--         --    for both Port A and Port B
--      c_use_ecc                => 0,
--         -- See DS512 for the limited core option selections for ECC support
--      c_use_ramb16bwer_rst_bhv => 0    --0, 1
--      )
--   port map
--      (
--      clka    => RX_CLIENT_CLK,
--      ssra    => RESET2RX_CLIENT,
--      dina    => rx_client_rxd_dpmem_wr_data_d1,
--      addra   => rx_client_rxd_dpmem_addr_d1,
--      ena     => rx_client_clk_enbl_d1,
--      regcea  => '0',
--      wea     => rx_client_rxd_dpmem_wr_en_d1,
--      douta   => RX_CLIENT_RXD_DPMEM_RD_DATA,
--
--
--      clkb    => AXI_STR_RXD_ACLK,
--      ssrb    => RESET2AXI_STR_RXD,
--      dinb    => AXI_STR_RXD_DPMEM_WR_DATA,
--      addrb   => AXI_STR_RXD_DPMEM_ADDR,
--      enb     => '1',
--      regceb  => '0',
--      web     => AXI_STR_RXD_DPMEM_WR_EN,
--      doutb   => AXI_STR_RXD_DPMEM_RD_DATA,
--
--      dbiterr => open,
--      sbiterr => open
--      );

I_RXS_MEM: xpm_memory_tdpram
  generic map (

    -- Common module generics
    MEMORY_SIZE             => 36*(C_RXS_MEM_BYTES/4),            --positive integer
    MEMORY_PRIMITIVE        => "block",          --string; "auto", "distributed", "block" or "ultra" ;
    CLOCKING_MODE           => "independent_clock",  --string; "common_clock", "independent_clock" 
    MEMORY_INIT_FILE        => "none",          --string; "none" or "<filename>.mem" 
    MEMORY_INIT_PARAM       => "",              --string;
    USE_MEM_INIT            => 1,               --integer; 0,1
    WAKEUP_TIME             => "disable_sleep", --string; "disable_sleep" or "use_sleep_pin" 
    MESSAGE_CONTROL         => 0,               --integer;
    ECC_MODE                => "no_ecc",        --string; "no_ecc", "encode_only", "decode_only" or "both_encode_and_decode" 
    AUTO_SLEEP_TIME         => 0,               --Do not Change
    USE_EMBEDDED_CONSTRAINT => 0,               --integer: 0,1
    MEMORY_OPTIMIZATION     => "true",          --string; "true", "false" 

    -- Port A module generics
    WRITE_DATA_WIDTH_A      => 36,              --positive integer
    READ_DATA_WIDTH_A       => 36,              --positive integer
    BYTE_WRITE_WIDTH_A      => 36,              --integer; 8, 9, or WRITE_DATA_WIDTH_A value
    ADDR_WIDTH_A            => (log2(C_RXS_MEM_BYTES/4)),               --positive integer
    READ_RESET_VALUE_A      => "0",             --string
    READ_LATENCY_A          => 1,               --non-negative integer
    WRITE_MODE_A            => "no_change",     --string; "write_first", "read_first", "no_change" 

    -- Port B module generics
    WRITE_DATA_WIDTH_B      => 36,              --positive integer
    READ_DATA_WIDTH_B       => 36,              --positive integer
    BYTE_WRITE_WIDTH_B      => 36,              --integer; 8, 9, or WRITE_DATA_WIDTH_B value
    ADDR_WIDTH_B            => (log2(C_RXS_MEM_BYTES/4)),               --positive integer
    READ_RESET_VALUE_B      => "0",             --string
    READ_LATENCY_B          => 1,               --non-negative integer
    WRITE_MODE_B            => "no_change"      --string; "write_first", "read_first", "no_change" 
  )
  port map (

    -- Common module ports
    sleep                   => '0',

    -- Port A module ports
    clka                    => RX_CLIENT_CLK,
    rsta                    => RESET2RX_CLIENT,
    ena                     => rx_client_clk_enbl_d1,
    regcea                  => '0',
    wea                     => rx_client_rxs_dpmem_wr_en_d1,
    addra                   => rx_client_rxs_dpmem_addr_d1,
    dina                    => rx_client_rxs_dpmem_wr_data_d1,
    injectsbiterra          => '0',
    injectdbiterra          => '0',
    douta                   => RX_CLIENT_RXS_DPMEM_RD_DATA,
    sbiterra                => open,
    dbiterra                => open,

    -- Port B module ports
    clkb                    => AXI_STR_RXS_ACLK,
    rstb                    => RESET2AXI_STR_RXS,
    enb                     => '1',
    regceb                  => '0',
    web                     => AXI_STR_RXS_DPMEM_WR_EN,
    addrb                   => AXI_STR_RXS_DPMEM_ADDR,
    dinb                    => AXI_STR_RXS_DPMEM_WR_DATA,
    injectsbiterrb          => '0',
    injectdbiterrb          => '0',
    doutb                   => AXI_STR_RXS_DPMEM_RD_DATA,
    sbiterrb                => open,
    dbiterrb                => open
  );

-- End of xpm_memory_tdpram_inst instance declaration

-- I_RXS_MEM : entity lib_bmg_v1_0.blk_mem_gen_wrapper
--   generic map(
--      c_family                 => C_FAMILY,
--      c_xdevicefamily          => C_FAMILY,
--
--      -- Selection between BMG and XPM
--      bmg_xpm_sel              => 0,
--      -- Memory Specific Configurations
--      c_mem_type               => 2,
--         -- This wrapper only supports the True Dual Port RAM
--         -- 0: Single Port RAM
--         -- 1: Simple Dual Port RAM
--         -- 2: True Dual Port RAM
--         -- 3: Single Port Rom
--         -- 4: Dual Port RAM
--      c_algorithm              => 1,
--         -- 0: Selectable Primative
--         -- 1: Minimum Area
--      c_prim_type              => 1,
--         -- 0: ( 1-bit wide)
--         -- 1: ( 2-bit wide)
--         -- 2: ( 4-bit wide)
--         -- 3: ( 9-bit wide)
--         -- 4: (18-bit wide)
--         -- 5: (36-bit wide)
--         -- 6: (72-bit wide, single port only)
--      c_byte_size              => 9,   -- 8 or 9
--
--      -- Simulation Behavior Options
--      c_sim_collision_check    => "NONE",
--         -- "None"
--         -- "Generate_X"
--         -- "All"
--         -- "Warnings_only"
--      c_common_clk             => 0,   -- 0, 1
--      c_disable_warn_bhv_coll  => 0,   -- 0, 1
--      c_disable_warn_bhv_range => 0,   -- 0, 1
--
--      -- Initialization Configuration Options
--      c_load_init_file         => 0,
--      c_init_file_name         => "none",
--      c_use_default_data       => 0,   -- 0, 1
--      c_default_data           => "0", -- "..."
--
--      -- Port A Specific Configurations
--      c_has_mem_output_regs_a  => 0,   -- 0, 1
--      c_has_mux_output_regs_a  => 0,   -- 0, 1
--      c_write_width_a          => 36,  -- 1 to 1152
--      c_read_width_a           => 36,  -- 1 to 1152
--      c_write_depth_a          => (C_RXS_MEM_BYTES/4),  -- 2 to 9011200
--      c_read_depth_a           => (C_RXS_MEM_BYTES/4),  -- 2 to 9011200
--      c_addra_width            => (log2(C_RXS_MEM_BYTES/4)),   -- 1 to 24
--      c_write_mode_a           => "NO_CHANGE",
--         -- "Write_First"
--         -- "Read_first"
--         -- "No_Change"
--      c_has_ena                => 1,   -- 0, 1
--      c_has_regcea             => 0,   -- 0, 1
--      c_has_ssra               => 0,   -- 0, 1
--      c_sinita_val             => "0", --"..."
--      c_use_byte_wea           => 0,   -- 0, 1
--      c_wea_width              => 1,   -- 1 to 128
--
--      -- Port B Specific Configurations
--      c_has_mem_output_regs_b  => 0,   -- 0, 1
--      c_has_mux_output_regs_b  => 0,   -- 0, 1
--      c_write_width_b          => 36,  -- 1 to 1152
--      c_read_width_b           => 36,  -- 1 to 1152
--      c_write_depth_b          => (C_RXS_MEM_BYTES/4),  -- 2 to 9011200
--      c_read_depth_b           => (C_RXS_MEM_BYTES/4),   -- 2 to 9011200
--      c_addrb_width            => (log2(C_RXS_MEM_BYTES/4)),   -- 1 to 24
--      c_write_mode_b           => "NO_CHANGE",
--         -- "Write_First"
--         -- "Read_first"
--         -- "No_Change"
--      c_has_enb                => 0,   -- 0, 1
--      c_has_regceb             => 0,   -- 0, 1
--      c_has_ssrb               => 0,   -- 0, 1
--      c_sinitb_val             => "0", -- "..."
--      c_use_byte_web           => 0,   -- 0, 1
--      c_web_width              => 1,   -- 1 to 128
--
--      -- Other Miscellaneous Configurations
--      c_mux_pipeline_stages    => 0,   -- 0, 1, 2, 3
--         -- The number of pipeline stages within the MUX
--         --    for both Port A and Port B
--      c_use_ecc                => 0,
--         -- See DS512 for the limited core option selections for ECC support
--      c_use_ramb16bwer_rst_bhv => 0    --0, 1
--      )
--   port map
--      (
--      clka    => RX_CLIENT_CLK,
--      ssra    => RESET2RX_CLIENT,
--      dina    => rx_client_rxs_dpmem_wr_data_d1,
--      addra   => rx_client_rxs_dpmem_addr_d1,
--      ena     => rx_client_clk_enbl_d1,
--      regcea  => '0',
--      wea     => rx_client_rxs_dpmem_wr_en_d1,
--      douta   => RX_CLIENT_RXS_DPMEM_RD_DATA,
--
--
--      clkb    => AXI_STR_RXS_ACLK,
--      ssrb    => RESET2AXI_STR_RXS,
--      dinb    => AXI_STR_RXS_DPMEM_WR_DATA,
--      addrb   => AXI_STR_RXS_DPMEM_ADDR,
--      enb     => '1',
--      regceb  => '0',
--      web     => AXI_STR_RXS_DPMEM_WR_EN,
--      doutb   => AXI_STR_RXS_DPMEM_RD_DATA,
--
--      dbiterr => open,
--      sbiterr => open
--      );

end rtl;


------------------------------------------------------------------------------
-- rx_if.vhd
------------------------------------------------------------------------------
--
-- *************************************************************************
--
-- (c) Copyright 2004-2011 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-- *************************************************************************
--
-- ------------------------------------------------------------------------------
--
------------------------------------------------------------------------------
-- Filename:        rx_if.vhd
-- Description:     Receive interface between AXIStream and Temac
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to rtlrove
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:          MSH
--
--  MSH     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of : out   std_logic; port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Libraries used;
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.rx_if_pack.all;

-------------------------------------------------------------------------------
-- Definition of Generics :
-------------------------------------------------------------------------------
-- System generics
--  C_FAMILY              -- Xilinx FPGA Family
--
-- Ethernet generics
--  C_HAS_SGMII
--     SGMII is the only PHY mode which causes a change in this Rx logic.
--  C_RXCSUM
--     0  No checksum offloading
--     1  Partial (legacy) checksum offloading
--     2  Full checksum offloading
--  C_RXVLAN_TRAN         -- Enable RX enhanced VLAN translation
--  C_RXVLAN_TAG          -- Enable RX enhanced VLAN taging
--  C_RXVLAN_STRP         -- Enable RX enhanced VLAN striping
--  C_MCAST_EXTEND        -- Enable RX extended multicast address filtering

-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Definition of Ports :
-------------------------------------------------------------------------------
--    BUS2IP_CLK
--    BUS2IP_RESET
--
--    AXI_STR_RXD_ACLK
--    AXI_STR_RXD_VALID
--    AXI_STR_RXD_READY
--    AXI_STR_RXD_LAST
--    AXI_STR_RXD_STRB
--    AXI_STR_RXD_DATA
--
--    AXI_STR_RXS_ACLK
--    AXI_STR_RXS_VALID
--    AXI_STR_RXS_READY
--    AXI_STR_RXS_LAST
--    AXI_STR_RXS_STRB
--    AXI_STR_RXS_DATA
--
--    EMAC_CLIENT_RXD_LEGACY
--    EMAC_CLIENT_RXD_VLD_LEGACY
--    EMAC_CLIENT_RX_GOODFRAME_LEGACY
--    EMAC_CLIENT_RX_BADFRAME_LEGACY
--    EMAC_CLIENT_RX_FRAMEDROP
--    LEGACY_RX_FILTER_MATCH
--
--    RX_CLIENT_CLK
--    RX_CLIENT_CLK_ENBL
--
--    EMAC_CLIENT_RX_STATS
--    EMAC_CLIENT_RX_STATS_VLD
--    EMAC_CLIENT_RX_STATS_BYTE_VLD
--    EMAC_CLIENT_RXD_VLD_2STATS
--    SOFT_EMAC_CLIENT_RX_STATS
--
--    RTAGREGDATA
--    TPID0REGDATA
--    TPID1REGDATA
--    UAWLREGDATA
--    UAWUREGDATA
--    RXCLCLKMCASTADDR
--    RXCLCLKMCASTEN
--    RXCLCLKMCASTRDDATA
--    LLINKCLKVLANADDR
--    LLINKCLKVLANRDDATA
--    LLINKCLKRXVLANBRAMENA
--
--    LLINKCLKEMULTIFLTRENBL
--    LLINKCLKNEWFNCENBL
--    LLINKCLKRXVSTRPMODE
--    LLINKCLKRXVTAGMODE
-------------------------------------------------------------------------------
----                  Entity Section
-------------------------------------------------------------------------------

entity rx_if is
  generic (
    C_FAMILY              : string                        := "virtex6";
    C_HAS_SGMII           : integer range 0 to 1          := 0;
    C_RXCSUM              : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_RXMEM               : integer                       := 4096;
    C_RXVLAN_TRAN         : integer range 0 to 1          := 0;
    C_RXVLAN_TAG          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP         : integer range 0 to 1          := 0;
    C_ENABLE_1588         : integer   := 0;
    C_MCAST_EXTEND        : integer range 0 to 1          := 0
    );

  port    (
    RX_FRAME_RECEIVED_INTRPT        : out std_logic;                          --  Frame received interrupt
    RX_FRAME_REJECTED_INTRPT        : out std_logic;                          --  Frame rejected interrupt
    RX_BUFFER_MEM_OVERFLOW_INTRPT   : out std_logic;                          --  Memory overflow interrupt

    AXI_STR_RXD_ACLK                : in  std_logic;                          --  AXI-Stream Receive Data Clock
    AXI_STR_RXD_VALID               : out std_logic;                          --  AXI-Stream Receive Data Valid
    AXI_STR_RXD_READY               : in  std_logic;                          --  AXI-Stream Receive Data Ready
    AXI_STR_RXD_LAST                : out std_logic;                          --  AXI-Stream Receive Data Last
    AXI_STR_RXD_STRB                : out std_logic_vector(3 downto 0);       --  AXI-Stream Receive Data Keep
    AXI_STR_RXD_DATA                : out std_logic_vector(31 downto 0);      --  AXI-Stream Receive Data Data
    RESET2AXI_STR_RXD               : in  std_logic;                          --  AXI-Stream Receive Data Reset

    AXI_STR_RXS_ACLK                : in  std_logic;                          --  AXI-Stream Receive Status Clock
    AXI_STR_RXS_VALID               : out std_logic;                          --  AXI-Stream Receive Status Valid
    AXI_STR_RXS_READY               : in  std_logic;                          --  AXI-Stream Receive Status Ready
    AXI_STR_RXS_LAST                : out std_logic;                          --  AXI-Stream Receive Status Last
    AXI_STR_RXS_STRB                : out std_logic_vector(3 downto 0);       --  AXI-Stream Receive Status Keep
    AXI_STR_RXS_DATA                : out std_logic_vector(31 downto 0);      --  AXI-Stream Receive Status Data
    RESET2AXI_STR_RXS               : in  std_logic;                          --  AXI-Stream Receive Status Reset

    -- added 05/5/2011
    RX_CLK_ENABLE_IN                : in std_logic;                           -- TEMAC clock domain enable

    rx_statistics_vector            : in  std_logic_vector(27 downto 0);      -- RX statistics from TEMAC
    rx_statistics_valid             : in  std_logic;                          -- Rx stats valid from TEMAC
    rxspeedis10100                  : in  std_logic;                          -- speed is 10/100 not 1000 indicator

    rx_mac_aclk                     : in  std_logic;                          -- Rx axistream clock from TEMAC
    rx_reset                        : in  std_logic;                          -- Rx axistream reset from TEMAC
    rx_axis_mac_tdata               : in  std_logic_vector(7 downto 0);       -- Rx axistream data from TEMAC
    rx_axis_mac_tvalid              : in  std_logic;                          -- Rx axistream valid from TEMAC
    rx_axis_mac_tlast               : in  std_logic;                          -- Rx axistream last from TEMAC
    rx_axis_mac_tuser               : in  std_logic;                          -- Rx axistream good/bad indicator from TEMAC

    RX_CL_CLK_RX_TAG_REG_DATA       : in  std_logic_vector(0 to 31);          --  Receive VLAN TAG
    RX_CL_CLK_TPID0_REG_DATA        : in  std_logic_vector(0 to 31);          --  Receive VLAN TPID 0
    RX_CL_CLK_TPID1_REG_DATA        : in  std_logic_vector(0 to 31);          --  Receive VLAN TPID 1
    RX_CL_CLK_UAWL_REG_DATA         : in  std_logic_vector(0 to 31);          --  Receive Unicast Address Word Lower
    RX_CL_CLK_UAWU_REG_DATA         : in  std_logic_vector(16 to 31);         --  Receive Unicast Address Word Upper

    RX_CL_CLK_MCAST_ADDR            : out std_logic_vector(0 to 14);          --  Receive Multicast Memory Address
    RX_CL_CLK_MCAST_EN              : out std_logic;                          --  Receive Multicast Memory Address Enable
    RX_CL_CLK_MCAST_RD_DATA         : in  std_logic_vector(0 to 0);           --  Receive Multicast Memory Address Read Data

    RX_CL_CLK_VLAN_ADDR             : out std_logic_vector(0 to 11);          --  Receive VLAN Memory Address
    RX_CL_CLK_VLAN_RD_DATA          : in  std_logic_vector(18 to 31);         --  Receive VLAN Memory Read Data
    RX_CL_CLK_VLAN_BRAM_EN_A        : out std_logic;                          --  Receive VLAN Memory Enable

    RX_CL_CLK_BAD_FRAME_ENBL        : in  std_logic;                          --  Receive Bad Frame Enable
    RX_CL_CLK_EMULTI_FLTR_ENBL      : in  std_logic;                          --  Receive Extended Multicast Address Filter Enable
    RX_CL_CLK_NEW_FNC_ENBL          : in  std_logic;                          --  Receive New Function Enable
    RX_CL_CLK_BRDCAST_REJ           : in  std_logic;                          --  Receive Broadcast Reject
    RX_CL_CLK_MULCAST_REJ           : in  std_logic;                          --  Receive Multicast Reject
    RX_CL_CLK_VSTRP_MODE            : in  std_logic_vector(0 to 1);           --  Receive VLAN Strip Mode
    RX_CL_CLK_VTAG_MODE             : in  std_logic_vector(0 to 1)            --  Receive VLAN TAG Mode

    );
end rx_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture rtl of rx_if is

function log2(x : natural) return integer is
  variable i  : integer := 0;
  variable val: integer := 1;
begin
  if x = 0 then return 0;
  else
    for j in 0 to 29 loop -- for loop for XST 
      if val >= x then null;
      else
        i := i+1;
        val := val*2;
      end if;
    end loop;
  -- synthesis translate_off
    assert val >= x
      report "Function log2 received argument larger" &
             " than its capability of 2^30. "
      severity failure;
  -- synthesis translate_on
    return i;
  end if;
end function log2;

------------------------------------------------------------------------------
-- Constant Declarations
------------------------------------------------------------------------------

constant C_RXD_MEM_BYTES      : integer := C_RXMEM;
constant C_RXD_MEM_ADDR_WIDTH : integer := (log2(C_RXD_MEM_BYTES/4))-1;
constant C_RXS_MEM_BYTES      : integer := (C_RXMEM/2);
constant C_RXS_MEM_ADDR_WIDTH : integer := (log2(C_RXS_MEM_BYTES/4))-1;
constant C_RXVLAN_WIDTH       : integer := (C_RXVLAN_TRAN*12) + C_RXVLAN_TAG + C_RXVLAN_STRP;

------------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------------
type type_end_of_frame_reset_array is array (1 to 18) of std_logic;
signal end_of_frame_reset_array : type_end_of_frame_reset_array;
signal end_of_frame_reset_array_in : std_logic;

type RECEIVE_DATA_VALID_GEN_SM_TYPE is (
       IDLE,
       RECEIVING_NOW
     );
signal receive_data_valid_gen_current_state : RECEIVE_DATA_VALID_GEN_SM_TYPE;
signal receive_data_valid_gen_next_state    : RECEIVE_DATA_VALID_GEN_SM_TYPE;

signal axi_str_rxd_dpmem_wr_data       : std_logic_vector(35 downto 0);
signal axi_str_rxd_dpmem_rd_data       : std_logic_vector(35 downto 0);
signal axi_str_rxd_dpmem_wr_en         : std_logic_vector(0 downto 0);
signal axi_str_rxd_dpmem_addr          : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);

signal axi_str_rxs_dpmem_wr_data       : std_logic_vector(35 downto 0);
signal axi_str_rxs_dpmem_rd_data       : std_logic_vector(35 downto 0);
signal axi_str_rxs_dpmem_wr_en         : std_logic_vector(0 downto 0);
signal axi_str_rxs_dpmem_addr          : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);

signal rx_client_rxd_dpmem_wr_data     : std_logic_vector(35 downto 0);
signal rx_client_rxd_dpmem_rd_data     : std_logic_vector(35 downto 0);
signal rx_client_rxd_dpmem_wr_en       : std_logic_vector(0 downto 0);
signal rx_client_rxd_dpmem_addr        : std_logic_vector(C_RXD_MEM_ADDR_WIDTH downto 0);

signal rx_client_rxs_dpmem_wr_data     : std_logic_vector(35 downto 0);
signal rx_client_rxs_dpmem_rd_data     : std_logic_vector(35 downto 0);
signal rx_client_rxs_dpmem_wr_en       : std_logic_vector(0 downto 0);
signal rx_client_rxs_dpmem_addr        : std_logic_vector(C_RXS_MEM_ADDR_WIDTH downto 0);
signal axi_str_rxd_mem_last_read_out_ptr_gray : std_logic_vector(35 downto 0);
signal axi_str_rxs_mem_last_read_out_ptr_gray : std_logic_vector(35 downto 0);

signal derived_rx_good_frame_i         : std_logic;
signal derived_rx_bad_frame_i          : std_logic;
signal derived_rx_good_frame_d1        : std_logic;
signal derived_rx_bad_frame_d1         : std_logic;
signal derived_rx_good_frame           : std_logic;
signal derived_rx_bad_frame            : std_logic;
signal derived_rxd_vld                 : std_logic;
signal derived_rx_clk_enbl             : std_logic;
signal derived_rx_clk_enbl_reg1        : std_logic;
signal derived_rx_clk_enbl_reg2        : std_logic;
signal derived_rx_clk_enbl_cmb         : std_logic;

signal rx_axis_mac_tdata_d1            : std_logic_vector(7 downto 0);
signal rx_axis_mac_tvalid_d1           : std_logic;
signal rx_axis_mac_tlast_d1            : std_logic;
signal rx_axis_mac_tlast_d2            : std_logic;
signal rx_axis_mac_tlast_d3            : std_logic;
signal rx_axis_mac_tlast_d4           : std_logic;

signal rx_axis_mac_tvalid_d2           : std_logic;
signal rx_axis_mac_tvalid_d3           : std_logic;
signal rx_tvalid_start        : std_logic;
signal rx_tvalid_end          : std_logic;
signal rx_tvalid              : std_logic;
signal rx_tvalid_d1           : std_logic;
signal rx_tvalid_d2           : std_logic;
signal rx_tvalid_d3           : std_logic;
signal rx_tvalid_d4           : std_logic;
signal no_stripping           : std_logic;
signal no_stripping_d1        : std_logic;
signal no_stripping_d2        : std_logic;
signal no_stripping_d3        : std_logic;
signal rx_statistics_vector_i : std_logic_vector(27 downto 0);
signal rx_statistics_valid_i  : std_logic;
signal end_of_frame_pulse     : std_logic;

begin

  end_of_frame_reset_array_in  <= end_of_frame_reset_array(12);

  PIPE_ENDOFFRAMERESET : process (rx_mac_aclk)
  begin
   if rising_edge(rx_mac_aclk) then
     if rx_reset = '1' then
       end_of_frame_reset_array <= (others => '0');
     else
       if (derived_rx_clk_enbl = '1') then
         end_of_frame_reset_array (1)  <= end_of_frame_pulse;
         for i in 1 to 17 loop
           end_of_frame_reset_array (i+1) <= end_of_frame_reset_array (i);
         end loop;
       end if;
     end if;
   end if;
  end process;

  -- Create end of frame reset using TLAST which does not move in relationship
  -- to the next frame coming in.

  ENDOFFRAMEPULSE_PROCESS : process (rx_mac_aclk)
  begin
   if rising_edge(rx_mac_aclk) then
     if rx_reset = '1' then
       end_of_frame_pulse <= '0';
     else
       end_of_frame_pulse <= rx_axis_mac_tlast or           -- set when tlast indicates end of frame
         (end_of_frame_pulse and                            -- hold until the next clock enable
         not (end_of_frame_pulse and derived_rx_clk_enbl)); -- clear next clock enable after set
     end if;
   end if;
  end process;

  -- capture statistics valid and statistics until end of frame reset because in
  -- MGT 10/100Mbps modes the clock enable does not exist when this comes out if
  -- fcs stripping is enabled and it is missed in the next level down
  CAPTURE_STATS_PROCESS : process(rx_mac_aclk)
  begin
   if rising_edge(rx_mac_aclk) then
     if rx_reset = '1' then
        rx_statistics_vector_i <= (others => '0');
        rx_statistics_valid_i  <= '0';
      else
        if (rx_axis_mac_tlast_d4 = '1') then
          rx_statistics_vector_i <= (others => '0');
          rx_statistics_valid_i  <= '0';
        elsif (rx_statistics_valid = '1') then
          rx_statistics_vector_i <= rx_statistics_vector;
          rx_statistics_valid_i  <= '1';
        else
          NULL;
        end if;
      end if;
    end if;
  end process CAPTURE_STATS_PROCESS;

  derived_rx_good_frame_i <= rx_axis_mac_tlast and not(rx_axis_mac_tuser);
  derived_rx_bad_frame_i  <= rx_axis_mac_tlast and    (rx_axis_mac_tuser);

   -- stretch good bad for 10/100 clock enable case
  STRETCH_GOOD_BAD_PROCESS : process(rx_mac_aclk)
  begin
   if rising_edge(rx_mac_aclk) then
     if rx_reset = '1' then
        derived_rx_good_frame_d1 <= '0';
        derived_rx_bad_frame_d1  <= '0';
      else
        derived_rx_good_frame_d1 <= derived_rx_good_frame_i;
        derived_rx_bad_frame_d1  <= derived_rx_bad_frame_i;
      end if;
    end if;
  end process STRETCH_GOOD_BAD_PROCESS;

  derived_rx_good_frame <= derived_rx_good_frame_i or derived_rx_good_frame_d1;
  derived_rx_bad_frame  <= derived_rx_bad_frame_i  or derived_rx_bad_frame_d1;

  --------------------------------------------------------------------------
  -- receive data valid gen State Machine
  -- RXDVLDSM_REGS_PROCESS: registered process of the state machine
  -- RXDVLDSM_CMB_PROCESS:  combinatorial next-state logic
  --------------------------------------------------------------------------

  RXDVLDSM_REGS_PROCESS: process (rx_mac_aclk)
  begin
    if rising_edge(rx_mac_aclk) then
      if rx_reset = '1' then
        receive_data_valid_gen_current_state <= IDLE;
        derived_rx_clk_enbl_reg1 <= '0';
        derived_rx_clk_enbl_reg2 <= '0';
      else
        receive_data_valid_gen_current_state <= receive_data_valid_gen_next_state;
        derived_rx_clk_enbl_reg1 <= derived_rx_clk_enbl_cmb after 1 ps;
        derived_rx_clk_enbl_reg2 <= derived_rx_clk_enbl_reg1 after 1 ps;
      end if;
    end if;
  end process;

  NOT_SGMII: if(C_HAS_SGMII = 0) generate
    derived_rx_clk_enbl <= '1' when rxspeedis10100 = '0' else -- speed is 1000
                           RX_CLK_ENABLE_IN;                                                                     -- speed is 10 or 100
  end generate NOT_SGMII;

  IS_SGMII: if(C_HAS_SGMII = 1) generate
    derived_rx_clk_enbl <= '1' when rxspeedis10100 = '0' else -- speed is 1000
                           derived_rx_clk_enbl_reg1;                                                             -- speed is 10 or 100
  end generate IS_SGMII;

  RXDVLDSM_CMB_PROCESS: process (
    RX_CLK_ENABLE_IN,
    rx_axis_mac_tvalid,
    rx_axis_mac_tlast,
    receive_data_valid_gen_current_state
    )
  begin

    case receive_data_valid_gen_current_state is

      when IDLE =>
        if (rx_axis_mac_tvalid = '1') then
          receive_data_valid_gen_next_state <= RECEIVING_NOW;
          derived_rx_clk_enbl_cmb           <= rx_axis_mac_tvalid;
        else
          receive_data_valid_gen_next_state <= IDLE;
          derived_rx_clk_enbl_cmb           <= RX_CLK_ENABLE_IN;
        end if;

      when RECEIVING_NOW =>
        if (rx_axis_mac_tlast = '1') then
          receive_data_valid_gen_next_state <= IDLE;
          derived_rx_clk_enbl_cmb           <= rx_axis_mac_tvalid;
        else
          receive_data_valid_gen_next_state <= RECEIVING_NOW;
          derived_rx_clk_enbl_cmb           <= rx_axis_mac_tvalid;
        end if;

      when others   =>
        receive_data_valid_gen_next_state   <= IDLE;
        derived_rx_clk_enbl_cmb             <= RX_CLK_ENABLE_IN;
    end case;
  end process;

  detect_stripping: process (rx_mac_aclk)
  begin
    if rising_edge(rx_mac_aclk) then
      if rx_reset = '1' then
        no_stripping    <= '0';
        no_stripping_d1 <= '0';
        no_stripping_d2 <= '0';
        no_stripping_d3 <= '0';
      elsif (rx_axis_mac_tlast = '1') and (rx_tvalid_d1 = '1') then
        no_stripping    <= '1';
        no_stripping_d1 <= no_stripping;
        no_stripping_d2 <= no_stripping_d1;
        no_stripping_d3 <= no_stripping_d2;
      elsif (rx_tvalid_end = '1' or rx_tvalid_d4 = '1') then
        no_stripping    <= '0';
        no_stripping_d1 <= no_stripping;
        no_stripping_d2 <= no_stripping_d1;
        no_stripping_d3 <= no_stripping_d2;
      else
        no_stripping    <= no_stripping;
        no_stripping_d1 <= no_stripping;
        no_stripping_d2 <= no_stripping_d1;
        no_stripping_d3 <= no_stripping_d2;
      end if;
    end if;
   end process detect_stripping;

  CREATE_RXD_VLD_PROCESS: process (rx_mac_aclk)
  begin
    if rising_edge(rx_mac_aclk) then
      if rx_reset = '1' then
        derived_rxd_vld       <= '0';
        rx_axis_mac_tdata_d1  <= (others => '0');
        rx_axis_mac_tvalid_d1 <= '0';
        rx_axis_mac_tvalid_d2    <= '0';
        rx_axis_mac_tvalid_d3    <= '0';
        rx_axis_mac_tlast_d1     <= '0';
        rx_axis_mac_tlast_d2     <= '0';
        rx_axis_mac_tlast_d3     <= '0';
        rx_axis_mac_tlast_d4     <= '0';
        rx_tvalid_start <= '0';
        rx_tvalid_end   <= '0';
        rx_tvalid       <= '0';
        rx_tvalid_d1    <= '0';
        rx_tvalid_d2    <= '0';
        rx_tvalid_d3    <= '0';
        rx_tvalid_d4    <= '0';
      else
        rx_tvalid_d1    <= rx_tvalid;
        rx_tvalid_d2    <= rx_tvalid_d1;
        rx_tvalid_d3    <= rx_tvalid_d2;
        rx_tvalid_d4    <= rx_tvalid_d3;

        if (rx_axis_mac_tvalid = '0') and (rx_axis_mac_tvalid_d1 = '0') and (rx_axis_mac_tvalid_d3 = '1') then
          rx_tvalid_end <= '1';
        else
          rx_tvalid_end <= '0';
        end if;

        if (rx_axis_mac_tvalid = '1') and (rx_axis_mac_tvalid_d1 = '0') and (rx_axis_mac_tvalid_d2 = '0') and
           (rx_axis_mac_tvalid_d3 = '0') and (rx_axis_mac_tlast = '0')then
          rx_tvalid_start <= '1';
        else
          rx_tvalid_start <= '0';
        end if;

        if rxspeedis10100 = '1' then -- speed is 10 or 100 clock enable toggles
          if ((rx_axis_mac_tvalid = '1') and (rx_axis_mac_tvalid_d1 = '0') and (rx_axis_mac_tvalid_d2 = '0') and
              (rx_axis_mac_tvalid_d3 = '0') and (rx_axis_mac_tlast = '0')) then
            rx_tvalid <= '1';
          elsif (rx_tvalid_end = '1') then
            rx_tvalid <= '0';
          else
            null;
          end if;

          if (C_HAS_SGMII = 0) then -- not SGMII at 10/100
            if no_stripping_d2 = '1' or no_stripping_d3 = '1' then --terminate early if no fcs stripping
              derived_rxd_vld  <= '0';
            else
              derived_rxd_vld  <= rx_tvalid; -- extend to cover last byte when fcs stripping
            end if;

            if (rx_axis_mac_tvalid_d1 = '1' or rx_axis_mac_tvalid_d3 = '1') then
              rx_axis_mac_tdata_d1  <= rx_axis_mac_tdata;
            end if;
          else -- is SGMII at 10/100
            if no_stripping_d2 = '1' or no_stripping_d3 = '1'  or rx_axis_mac_tlast_d1 = '1' then --terminate early if no fcs strip
              derived_rxd_vld  <= '0';
            elsif (rx_axis_mac_tvalid = '1') then
              derived_rxd_vld  <= '1';
            else
              NULL;
            end if;

            rx_axis_mac_tdata_d1  <= rx_axis_mac_tdata;
          end if;

        else -- speed is 1000 clock enable always 1
          if rx_axis_mac_tlast = '1' and rx_axis_mac_tvalid_d1 = '0' then
            derived_rxd_vld  <= '0';
          else
            derived_rxd_vld  <= rx_axis_mac_tvalid or rx_axis_mac_tvalid_d1;
          end if;

          rx_axis_mac_tdata_d1  <= rx_axis_mac_tdata;
        end if;

        rx_axis_mac_tlast_d1     <= rx_axis_mac_tlast;
        rx_axis_mac_tlast_d2     <= rx_axis_mac_tlast_d1;
        rx_axis_mac_tlast_d3     <= rx_axis_mac_tlast_d2;
        rx_axis_mac_tlast_d4     <= rx_axis_mac_tlast_d3;

        if rx_axis_mac_tlast = '1' then
          rx_axis_mac_tvalid_d1 <= '0';
          rx_axis_mac_tvalid_d2 <= rx_axis_mac_tvalid_d1;
          rx_axis_mac_tvalid_d3 <= rx_axis_mac_tvalid_d2;
        else
          rx_axis_mac_tvalid_d1 <= rx_axis_mac_tvalid;
          rx_axis_mac_tvalid_d2 <= rx_axis_mac_tvalid_d1;
          rx_axis_mac_tvalid_d3 <= rx_axis_mac_tvalid_d2;
        end if;
      end if;
    end if;
  end process CREATE_RXD_VLD_PROCESS;
  RX_DP_MEM_IF_I : rx_mem_if
  generic map (
    C_RXD_MEM_BYTES      => C_RXD_MEM_BYTES,
    C_RXD_MEM_ADDR_WIDTH => C_RXD_MEM_ADDR_WIDTH,
    C_RXS_MEM_BYTES      => C_RXS_MEM_BYTES,
    C_RXS_MEM_ADDR_WIDTH => C_RXS_MEM_ADDR_WIDTH,
    C_FAMILY             => C_FAMILY
  )
  port map(
    AXI_STR_RXD_ACLK            => AXI_STR_RXD_ACLK,
    AXI_STR_RXD_DPMEM_WR_DATA   => axi_str_rxd_dpmem_wr_data,
    AXI_STR_RXD_DPMEM_RD_DATA   => axi_str_rxd_dpmem_rd_data,
    AXI_STR_RXD_DPMEM_WR_EN     => axi_str_rxd_dpmem_wr_en,
    AXI_STR_RXD_DPMEM_ADDR      => axi_str_rxd_dpmem_addr,
    RESET2AXI_STR_RXD           => RESET2AXI_STR_RXD,

    AXI_STR_RXS_ACLK            => AXI_STR_RXS_ACLK,
    AXI_STR_RXS_DPMEM_WR_DATA   => axi_str_rxs_dpmem_wr_data,
    AXI_STR_RXS_DPMEM_RD_DATA   => axi_str_rxs_dpmem_rd_data,
    AXI_STR_RXS_DPMEM_WR_EN     => axi_str_rxs_dpmem_wr_en,
    AXI_STR_RXS_DPMEM_ADDR      => axi_str_rxs_dpmem_addr,
    RESET2AXI_STR_RXS           => RESET2AXI_STR_RXS,

    RX_CLIENT_CLK               => rx_mac_aclk,
    RX_CLIENT_CLK_ENBL          => derived_rx_clk_enbl,
    RX_CLIENT_RXD_DPMEM_WR_DATA => rx_client_rxd_dpmem_wr_data,
    RX_CLIENT_RXD_DPMEM_RD_DATA => rx_client_rxd_dpmem_rd_data,
    RX_CLIENT_RXD_DPMEM_WR_EN   => rx_client_rxd_dpmem_wr_en,
    RX_CLIENT_RXD_DPMEM_ADDR    => rx_client_rxd_dpmem_addr,

    RX_CLIENT_RXS_DPMEM_WR_DATA => rx_client_rxs_dpmem_wr_data,
    RX_CLIENT_RXS_DPMEM_RD_DATA => rx_client_rxs_dpmem_rd_data,
    RX_CLIENT_RXS_DPMEM_WR_EN   => rx_client_rxs_dpmem_wr_en,
    RX_CLIENT_RXS_DPMEM_ADDR    => rx_client_rxs_dpmem_addr,
    RESET2RX_CLIENT         => rx_reset
  );

  NO_INCLUDE_RX_VLAN: if(C_RXVLAN_TRAN = 0 and C_RXVLAN_TAG = 0 and C_RXVLAN_STRP = 0) generate
  begin
    RX_EMAC_IF_I : rx_emac_if
    generic map (
      C_RXVLAN_WIDTH        => C_RXVLAN_WIDTH,
      C_RXD_MEM_BYTES       => C_RXD_MEM_BYTES,
      C_RXD_MEM_ADDR_WIDTH  => C_RXD_MEM_ADDR_WIDTH,
      C_RXS_MEM_BYTES       => C_RXS_MEM_BYTES,
      C_RXS_MEM_ADDR_WIDTH  => C_RXS_MEM_ADDR_WIDTH,
      C_FAMILY              => C_FAMILY,
      C_RXCSUM              => C_RXCSUM,
      C_RXVLAN_TRAN         => C_RXVLAN_TRAN,
      C_RXVLAN_TAG          => C_RXVLAN_TAG,
      C_RXVLAN_STRP         => C_RXVLAN_STRP,
      C_ENABLE_1588         => C_ENABLE_1588,
      C_MCAST_EXTEND        => C_MCAST_EXTEND
    )
    port map(
      RX_FRAME_RECEIVED_INTRPT        => RX_FRAME_RECEIVED_INTRPT,
      RX_FRAME_REJECTED_INTRPT        => RX_FRAME_REJECTED_INTRPT,
      RX_BUFFER_MEM_OVERFLOW_INTRPT   => RX_BUFFER_MEM_OVERFLOW_INTRPT,

      rx_statistics_vector            => rx_statistics_vector_i,
      rx_statistics_valid             => rx_statistics_valid_i,
      end_of_frame_reset_in           => end_of_frame_reset_array_in,

      rx_mac_aclk                     =>  rx_mac_aclk,
      rx_reset                        =>  rx_reset,
      derived_rxd                     =>  rx_axis_mac_tdata_d1,

      derived_rx_good_frame           =>  derived_rx_good_frame,
      derived_rx_bad_frame            =>  derived_rx_bad_frame,
      derived_rxd_vld                 =>  derived_rxd_vld,
      derived_rx_clk_enbl             =>  derived_rx_clk_enbl,

      RX_CL_CLK_RX_TAG_REG_DATA       => RX_CL_CLK_RX_TAG_REG_DATA,
      RX_CL_CLK_TPID0_REG_DATA        => RX_CL_CLK_TPID0_REG_DATA,
      RX_CL_CLK_TPID1_REG_DATA        => RX_CL_CLK_TPID1_REG_DATA,
      RX_CL_CLK_UAWL_REG_DATA         => RX_CL_CLK_UAWL_REG_DATA,
      RX_CL_CLK_UAWU_REG_DATA         => RX_CL_CLK_UAWU_REG_DATA,

      RX_CL_CLK_MCAST_ADDR            => RX_CL_CLK_MCAST_ADDR,
      RX_CL_CLK_MCAST_EN              => RX_CL_CLK_MCAST_EN,
      RX_CL_CLK_MCAST_RD_DATA         => RX_CL_CLK_MCAST_RD_DATA,

      RX_CL_CLK_VLAN_ADDR             => RX_CL_CLK_VLAN_ADDR,
      RX_CL_CLK_VLAN_RD_DATA          => RX_CL_CLK_VLAN_RD_DATA,
      RX_CL_CLK_VLAN_BRAM_EN_A        => RX_CL_CLK_VLAN_BRAM_EN_A,

      RX_CL_CLK_BAD_FRAME_ENBL        => RX_CL_CLK_BAD_FRAME_ENBL,
      RX_CL_CLK_EMULTI_FLTR_ENBL      => RX_CL_CLK_EMULTI_FLTR_ENBL,
      RX_CL_CLK_NEW_FNC_ENBL          => RX_CL_CLK_NEW_FNC_ENBL,
      RX_CL_CLK_BRDCAST_REJ           => RX_CL_CLK_BRDCAST_REJ,
      RX_CL_CLK_MULCAST_REJ           => RX_CL_CLK_MULCAST_REJ,
      RX_CL_CLK_VSTRP_MODE            => RX_CL_CLK_VSTRP_MODE,
      RX_CL_CLK_VTAG_MODE             => RX_CL_CLK_VTAG_MODE,

      RX_CLIENT_RXD_DPMEM_WR_DATA     => rx_client_rxd_dpmem_wr_data,
      RX_CLIENT_RXD_DPMEM_RD_DATA     => rx_client_rxd_dpmem_rd_data,
      RX_CLIENT_RXD_DPMEM_WR_EN       => rx_client_rxd_dpmem_wr_en,
      RX_CLIENT_RXD_DPMEM_ADDR        => rx_client_rxd_dpmem_addr,
      RX_CLIENT_RXS_DPMEM_WR_DATA     => rx_client_rxs_dpmem_wr_data,
      RX_CLIENT_RXS_DPMEM_RD_DATA     => rx_client_rxs_dpmem_rd_data,
      RX_CLIENT_RXS_DPMEM_WR_EN       => rx_client_rxs_dpmem_wr_en,
      RX_CLIENT_RXS_DPMEM_ADDR        => rx_client_rxs_dpmem_addr,

      AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY => axi_str_rxs_mem_last_read_out_ptr_gray,
      AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY => axi_str_rxd_mem_last_read_out_ptr_gray
    );
  end generate NO_INCLUDE_RX_VLAN;

  INCLUDE_RX_VLAN: if(C_RXVLAN_TRAN = 1 or C_RXVLAN_TAG = 1 or C_RXVLAN_STRP = 1) generate
  begin
    RX_EMAC_IF_I : rx_emac_if_vlan
    generic map (
      C_RXVLAN_WIDTH        => C_RXVLAN_WIDTH,
      C_RXD_MEM_BYTES       => C_RXD_MEM_BYTES,
      C_RXD_MEM_ADDR_WIDTH  => C_RXD_MEM_ADDR_WIDTH,
      C_RXS_MEM_BYTES       => C_RXS_MEM_BYTES,
      C_RXS_MEM_ADDR_WIDTH  => C_RXS_MEM_ADDR_WIDTH,
      C_FAMILY              => C_FAMILY,
      C_RXCSUM              => C_RXCSUM,
      C_RXVLAN_TRAN         => C_RXVLAN_TRAN,
      C_RXVLAN_TAG          => C_RXVLAN_TAG,
      C_RXVLAN_STRP         => C_RXVLAN_STRP,
      C_MCAST_EXTEND        => C_MCAST_EXTEND
    )
    port map(
      RX_FRAME_RECEIVED_INTRPT        => RX_FRAME_RECEIVED_INTRPT,
      RX_FRAME_REJECTED_INTRPT        => RX_FRAME_REJECTED_INTRPT,
      RX_BUFFER_MEM_OVERFLOW_INTRPT   => RX_BUFFER_MEM_OVERFLOW_INTRPT,

      rx_statistics_vector            => rx_statistics_vector_i,
      rx_statistics_valid             => rx_statistics_valid_i,
      end_of_frame_reset_in           => end_of_frame_reset_array_in,

      rx_mac_aclk                     =>  rx_mac_aclk,
      rx_reset                        =>  rx_reset,
      derived_rxd                     =>  rx_axis_mac_tdata_d1,

      derived_rx_good_frame           =>  derived_rx_good_frame,
      derived_rx_bad_frame            =>  derived_rx_bad_frame,
      derived_rxd_vld                 =>  derived_rxd_vld,
      derived_rx_clk_enbl             =>  derived_rx_clk_enbl,

      RX_CL_CLK_RX_TAG_REG_DATA       => RX_CL_CLK_RX_TAG_REG_DATA,
      RX_CL_CLK_TPID0_REG_DATA        => RX_CL_CLK_TPID0_REG_DATA,
      RX_CL_CLK_TPID1_REG_DATA        => RX_CL_CLK_TPID1_REG_DATA,
      RX_CL_CLK_UAWL_REG_DATA         => RX_CL_CLK_UAWL_REG_DATA,
      RX_CL_CLK_UAWU_REG_DATA         => RX_CL_CLK_UAWU_REG_DATA,

      RX_CL_CLK_MCAST_ADDR            => RX_CL_CLK_MCAST_ADDR,
      RX_CL_CLK_MCAST_EN              => RX_CL_CLK_MCAST_EN,
      RX_CL_CLK_MCAST_RD_DATA         => RX_CL_CLK_MCAST_RD_DATA,

      RX_CL_CLK_VLAN_ADDR             => RX_CL_CLK_VLAN_ADDR,
      RX_CL_CLK_VLAN_RD_DATA          => RX_CL_CLK_VLAN_RD_DATA,
      RX_CL_CLK_VLAN_BRAM_EN_A        => RX_CL_CLK_VLAN_BRAM_EN_A,

      RX_CL_CLK_BAD_FRAME_ENBL        => RX_CL_CLK_BAD_FRAME_ENBL,
      RX_CL_CLK_EMULTI_FLTR_ENBL      => RX_CL_CLK_EMULTI_FLTR_ENBL,
      RX_CL_CLK_NEW_FNC_ENBL          => RX_CL_CLK_NEW_FNC_ENBL,
      RX_CL_CLK_BRDCAST_REJ           => RX_CL_CLK_BRDCAST_REJ,
      RX_CL_CLK_MULCAST_REJ           => RX_CL_CLK_MULCAST_REJ,
      RX_CL_CLK_VSTRP_MODE            => RX_CL_CLK_VSTRP_MODE,
      RX_CL_CLK_VTAG_MODE             => RX_CL_CLK_VTAG_MODE,

      RX_CLIENT_RXD_DPMEM_WR_DATA     => rx_client_rxd_dpmem_wr_data,
      RX_CLIENT_RXD_DPMEM_RD_DATA     => rx_client_rxd_dpmem_rd_data,
      RX_CLIENT_RXD_DPMEM_WR_EN       => rx_client_rxd_dpmem_wr_en,
      RX_CLIENT_RXD_DPMEM_ADDR        => rx_client_rxd_dpmem_addr,
      RX_CLIENT_RXS_DPMEM_WR_DATA     => rx_client_rxs_dpmem_wr_data,
      RX_CLIENT_RXS_DPMEM_RD_DATA     => rx_client_rxs_dpmem_rd_data,
      RX_CLIENT_RXS_DPMEM_WR_EN       => rx_client_rxs_dpmem_wr_en,
      RX_CLIENT_RXS_DPMEM_ADDR        => rx_client_rxs_dpmem_addr,

      AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY => axi_str_rxs_mem_last_read_out_ptr_gray,
      AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY => axi_str_rxd_mem_last_read_out_ptr_gray
    );
  end generate INCLUDE_RX_VLAN;

  RX_AXISTREAM_IF_I : rx_axistream_if
  generic map (
    C_RXD_MEM_BYTES      => C_RXD_MEM_BYTES,
    C_RXD_MEM_ADDR_WIDTH => C_RXD_MEM_ADDR_WIDTH,
    C_RXS_MEM_BYTES      => C_RXS_MEM_BYTES,
    C_RXS_MEM_ADDR_WIDTH => C_RXS_MEM_ADDR_WIDTH,
    C_FAMILY             => C_FAMILY,
    C_RXCSUM             => C_RXCSUM,
    C_RXVLAN_TRAN        => C_RXVLAN_TRAN,
    C_RXVLAN_TAG         => C_RXVLAN_TAG,
    C_RXVLAN_STRP        => C_RXVLAN_STRP,
    C_MCAST_EXTEND       => C_MCAST_EXTEND
  )
  port map(
    AXI_STR_RXD_ACLK                => AXI_STR_RXD_ACLK,
    AXI_STR_RXD_VALID               => AXI_STR_RXD_VALID,
    AXI_STR_RXD_READY               => AXI_STR_RXD_READY,
    AXI_STR_RXD_LAST                => AXI_STR_RXD_LAST,
    AXI_STR_RXD_STRB                => AXI_STR_RXD_STRB,
    AXI_STR_RXD_DATA                => AXI_STR_RXD_DATA,
    RESET2AXI_STR_RXD               => RESET2AXI_STR_RXD,

    AXI_STR_RXS_ACLK                => AXI_STR_RXS_ACLK,
    AXI_STR_RXS_VALID               => AXI_STR_RXS_VALID,
    AXI_STR_RXS_READY               => AXI_STR_RXS_READY,
    AXI_STR_RXS_LAST                => AXI_STR_RXS_LAST,
    AXI_STR_RXS_STRB                => AXI_STR_RXS_STRB,
    AXI_STR_RXS_DATA                => AXI_STR_RXS_DATA,
    RESET2AXI_STR_RXS               => RESET2AXI_STR_RXS,

    AXI_STR_RXD_DPMEM_WR_DATA       => axi_str_rxd_dpmem_wr_data,
    AXI_STR_RXD_DPMEM_RD_DATA       => axi_str_rxd_dpmem_rd_data,
    AXI_STR_RXD_DPMEM_WR_EN         => axi_str_rxd_dpmem_wr_en,
    AXI_STR_RXD_DPMEM_ADDR          => axi_str_rxd_dpmem_addr,

    AXI_STR_RXS_DPMEM_WR_DATA       => axi_str_rxs_dpmem_wr_data,
    AXI_STR_RXS_DPMEM_RD_DATA       => axi_str_rxs_dpmem_rd_data,
    AXI_STR_RXS_DPMEM_WR_EN         => axi_str_rxs_dpmem_wr_en,
    AXI_STR_RXS_DPMEM_ADDR          => axi_str_rxs_dpmem_addr,

      AXI_STR_RXS_MEM_LAST_READ_OUT_PTR_GRAY => axi_str_rxs_mem_last_read_out_ptr_gray,
    AXI_STR_RXD_MEM_LAST_READ_OUT_PTR_GRAY => axi_str_rxd_mem_last_read_out_ptr_gray
  );

end rtl;


-------------------------------------------------------------------------------
-- tx_if - entity/architecture pair
-------------------------------------------------------------------------------
--
-- (c) Copyright 2010 - 2010 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-------------------------------------------------------------------------------
-- Filename:        tx_if.vhd
-- Version:         v1.00a
-- Description:     top level of embedded ip AXI Stream Transmit interface
--
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   This section shows the hierarchical structure of axi_ethernet.
--
--              axi_ethernet.vhd
--                axi_ethernt_soft_temac_wrap.vhd
--                axi_lite_ipif.vhd
--                embedded_top.vhd
--          ->      tx_if.vhd
--                    tx_axistream_if.vhd
--                    tx_mem_if
--                    tx_emac_if.vhd
--
-------------------------------------------------------------------------------
-- Author:          MW
--
--  MW     07/01/10
-- ^^^^^^
--  - Initial release of v1.00.a
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

library work;
use work.tx_if_pack.all;

-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity tx_if is
  generic (
    C_FAMILY               : string                        := "virtex6";
    C_HALFDUP              : integer range 0 to 1          := 0;
    C_TXCSUM               : integer range 0 to 2          := 0;
    C_TXMEM                : integer                       := 4096;
    C_ENABLE_1588          : integer   := 0;
    C_TXVLAN_TRAN          : integer range 0 to 1          := 0;
    C_SPEED_2P5            : integer range 0 to 1          := 0;
    C_TXVLAN_TAG           : integer range 0 to 1          := 0;
    C_TXVLAN_STRP          : integer range 0 to 1          := 0;
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32        := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32        := 32
  );
  port (

    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK                 : in  std_logic;                                     --  AXI-Stream Transmit Data Clk
    reset2axi_str_txd                : in  std_logic;                                     --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID               : in  std_logic;                                     --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY               : out std_logic;                                     --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST                : in  std_logic;                                     --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TSTRB                : in  std_logic_vector(3 downto 0);                  --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA                : in  std_logic_vector(31 downto 0);                 --  AXI-Stream Transmit Data Data
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK                 : in  std_logic;                                     --  AXI-Stream Transmit Control Clk
    reset2axi_str_txc                : in  std_logic;                                     --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID               : in  std_logic;                                     --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY               : out std_logic;                                     --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST                : in  std_logic;                                     --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TSTRB                : in  std_logic_vector(3 downto 0);                  --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA                : in  std_logic_vector(31 downto 0);                 --  AXI-Stream Transmit Control Data

    -- VLAN Interface
    tx_vlan_bram_addr                : out std_logic_vector(11 downto 0);                 --  Transmit VLAN BRAM Addr
    tx_vlan_bram_din                 : in  std_logic_vector(13 downto 0);                 --  Transmit VLAN BRAM Rd Data
    tx_vlan_bram_en                  : out std_logic;                                     --  Transmit VLAN BRAM Enable

    enable_newFncEn                  : out std_logic; --Only perform VLAN when FLAG = 0xA --  Enable Extended VLAN Functions
    transMode_cross                  : in  std_logic;                                     --  VLAN Translation Mode Control Bit
    tagMode_cross                    : in  std_logic_vector( 1 downto 0);                 --  VLAN TAG Mode Control Bits
    strpMode_cross                   : in  std_logic_vector( 1 downto 0);                 --  VLAN Strip Mode Control Bits

    tpid0_cross                      : in  std_logic_vector(15 downto 0);                 --  VLAN TPID
    tpid1_cross                      : in  std_logic_vector(15 downto 0);                 --  VLAN TPID
    tpid2_cross                      : in  std_logic_vector(15 downto 0);                 --  VLAN TPID
    tpid3_cross                      : in  std_logic_vector(15 downto 0);                 --  VLAN TPID

    newTagData_cross                 : in  std_logic_vector(31 downto 0);                 --  VLAN Tag Data

    tx_init_in_prog                  : out std_logic;                                     --  Tx is Initializing after a reset
    tx_init_in_prog_cross            : in  std_logic;                                     --  Tx is Initializing after a reset



    tx_mac_aclk                      : in  std_logic;                                 --  Tx AXI-Stream clock in
    tx_reset                         : in  std_logic;                                 --  take to reset combiner
    tx_axis_mac_tdata                : out std_logic_vector(7 downto 0);              --  Tx AXI-Stream data
    tx_axis_mac_tvalid               : out std_logic;                                 --  Tx AXI-Stream valid
    tx_axis_mac_tlast                : out std_logic;                                 --  Tx AXI-Stream last
    tx_axis_mac_tuser                : out std_logic;                  -- this is always driven low since an underflow cannot occur
    tx_axis_mac_tready               : in  std_logic;                                 --  Tx AXI-Stream ready in from TEMAC
    tx_collision                     : in  std_logic;                                 --  collision not used
    tx_retransmit                    : in  std_logic;                                 -- retransmit not used

    tx_client_10_100                 : in  std_logic;                                 --  Tx Client CE Toggles Indicator
    tx_cmplt                         : out std_logic                                  -- transmit is complete indicator

  );

end tx_if;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture imp of tx_if is

function log2(x : natural) return integer is
  variable i  : integer := 0;
  variable val: integer := 1;
begin
  if x = 0 then return 0;
  else
    for j in 0 to 29 loop -- for loop for XST 
      if val >= x then null;
      else
        i := i+1;
        val := val*2;
      end if;
    end loop;
  -- synthesis translate_off
    assert val >= x
      report "Function log2 received argument larger" &
             " than its capability of 2^30. "
      severity failure;
  -- synthesis translate_on
    return i;
  end if;
end function log2;

  signal tx_axis_mac_tdata_int   : std_logic_vector(7 downto 0);
  signal tx_axis_mac_tvalid_int  : std_logic;
  signal tx_axis_mac_tlast_int   : std_logic;
  signal tx_axis_mac_tuser_int   : std_logic;
  signal tx_axis_mac_tready_int  : std_logic;

  -- Read Port - AXI Stream Data
  constant c_TxD_write_width_a     : integer range  0 to 18       := (C_S_AXI_DATA_WIDTH + 4)/4;
  constant c_TxD_read_width_a      : integer range  0 to 18       := (C_S_AXI_DATA_WIDTH + 4)/4;
  constant c_TxD_write_depth_a     : integer range  0 to 32768    := C_TXMEM;
  constant c_TxD_read_depth_a      : integer range  0 to 32768    := C_TXMEM;
  constant c_TxD_addra_width       : integer range  0 to 15       := log2(C_TXMEM);
  constant c_TxD_wea_width         : integer range  0 to 2        := 1;
  --Write Port - AXI Stream Data
  constant c_TxD_write_width_b     : integer range 36 to 36       := C_S_AXI_DATA_WIDTH + 4;
  constant c_TxD_read_width_b      : integer range 36 to 36       := C_S_AXI_DATA_WIDTH + 4;
  constant c_TxD_write_depth_b     : integer range  0 to 8192     := C_TXMEM/4;
  constant c_TxD_read_depth_b      : integer range  0 to 8192     := C_TXMEM/4;
  constant c_TxD_addrb_width       : integer range  0 to 13       := log2(C_TXMEM/4);
  constant c_TxD_web_width         : integer range  0 to 4        := 4;

  --Read Port - AXI Stream Data
  signal Tx_Client_TxD_2_Mem_Din   : std_logic_vector(c_TxD_write_width_a -1 downto 0);
  signal Tx_Client_TxD_2_Mem_Addr  : std_logic_vector(c_TxD_addra_width   -1 downto 0);
  signal Tx_Client_TxD_2_Mem_Dout  : std_logic_vector(c_TxD_read_width_a  -1 downto 0);
  signal Tx_Client_TxD_2_Mem_En    : std_logic;
  signal Tx_Client_TxD_2_Mem_We    : std_logic_vector(c_TxD_wea_width     -1 downto 0);
  --Write Port - AXI Stream Data
  signal Axi_Str_TxD_2_Mem_Din     : std_logic_vector(c_TxD_write_width_b -1 downto 0);
  signal Axi_Str_TxD_2_Mem_Addr    : std_logic_vector(c_TxD_addrb_width   -1 downto 0);
  signal Axi_Str_TxD_2_Mem_Dout    : std_logic_vector(c_TxD_read_width_b  -1 downto 0);
  signal Axi_Str_TxD_2_Mem_En      : std_logic;
  signal Axi_Str_TxD_2_Mem_We      : std_logic_vector(c_TxD_web_width     -1 downto 0);

  --  Force to use only 1 BRAM for the device families
    --  V6 = 36K (36 x 1024)

  -- Read Port - AXI Stream Control
  constant c_TxC_write_width_a     : integer range 36 to 36       := C_S_AXI_DATA_WIDTH + 4;
  constant c_TxC_read_width_a      : integer range 36 to 36       := C_S_AXI_DATA_WIDTH + 4;
  constant c_TxC_write_depth_a     : integer range  0 to 1024     := 1024;
  constant c_TxC_read_depth_a      : integer range  0 to 1024     := 1024;
  constant c_TxC_addra_width       : integer range  0 to 10       := 10;
  constant c_TxC_wea_width         : integer range  0 to 1        := 1;
  --Write Port - AXI Stream Control
  constant c_TxC_write_width_b     : integer range 36 to 36       := C_S_AXI_DATA_WIDTH + 4;
  constant c_TxC_read_width_b      : integer range 36 to 36       := C_S_AXI_DATA_WIDTH + 4;
  constant c_TxC_write_depth_b     : integer range  0 to 1024     := 1024;
  constant c_TxC_read_depth_b      : integer range  0 to 1024     := 1024;
  constant c_TxC_addrb_width       : integer range  0 to 10       := 10;
  constant c_TxC_web_width         : integer range  0 to 1        := 1;

  --Read Port - AXI Stream Control
  signal Tx_Client_TxC_2_Mem_Din   : std_logic_vector(c_TxC_write_width_a -1 downto 0);
  signal Tx_Client_TxC_2_Mem_Addr  : std_logic_vector(c_TxC_addra_width   -1 downto 0);
  signal Tx_Client_TxC_2_Mem_Dout  : std_logic_vector(c_TxC_read_width_a  -1 downto 0);
  signal Tx_Client_TxC_2_Mem_En    : std_logic;
  signal Tx_Client_TxC_2_Mem_We    : std_logic_vector(c_TxC_wea_width     -1 downto 0);
  --Write Port - AXI Stream Control
  signal Axi_Str_TxC_2_Mem_Din     : std_logic_vector(c_TxC_write_width_b -1 downto 0);
  signal Axi_Str_TxC_2_Mem_Addr    : std_logic_vector(c_TxC_addrb_width   -1 downto 0);
  signal Axi_Str_TxC_2_Mem_Dout    : std_logic_vector(c_TxC_read_width_b  -1 downto 0);
  signal Axi_Str_TxC_2_Mem_En      : std_logic;
  signal Axi_Str_TxC_2_Mem_We      : std_logic_vector(c_TxC_web_width     -1 downto 0);


begin


        TX_AXISTREAM_INTERFACE : tx_axistream_if
        --  Interface for Transmit AxiStream Data and Control; and Tx Memory
        generic map (
          C_FAMILY               => C_FAMILY,
          C_HALFDUP              => C_HALFDUP,
          C_TXCSUM               => C_TXCSUM,
          C_TXMEM                => C_TXMEM,
          C_TXVLAN_TRAN          => C_TXVLAN_TRAN,
          C_TXVLAN_TAG           => C_TXVLAN_TAG,
          C_TXVLAN_STRP          => C_TXVLAN_STRP,
          C_S_AXI_ADDR_WIDTH     => C_S_AXI_ADDR_WIDTH,
          C_S_AXI_DATA_WIDTH     => C_S_AXI_DATA_WIDTH,

          -- Write Port - AXI Stream TxData
          c_TxD_write_width_b    => c_TxD_write_width_b,
          c_TxD_read_width_b     => c_TxD_read_width_b,
          c_TxD_write_depth_b    => c_TxD_write_depth_b,
          c_TxD_read_depth_b     => c_TxD_read_depth_b,
          c_TxD_addrb_width      => c_TxD_addrb_width,
          c_TxD_web_width        => c_TxD_web_width,

          -- Write Port - AXI Stream TxControl
          c_TxC_write_width_b    => c_TxC_write_width_b,
          c_TxC_read_width_b     => c_TxC_read_width_b,
          c_TxC_write_depth_b    => c_TxC_write_depth_b,
          c_TxC_read_depth_b     => c_TxC_read_depth_b,
          c_TxC_addrb_width      => c_TxC_addrb_width,
          c_TxC_web_width        => c_TxC_web_width

        )
        port map  (
          -- AXI Stream Data signals
          AXI_STR_TXD_ACLK       => AXI_STR_TXD_ACLK,
          reset2axi_str_txd      => reset2axi_str_txd,
          AXI_STR_TXD_TVALID     => AXI_STR_TXD_TVALID,
          AXI_STR_TXD_TREADY     => AXI_STR_TXD_TREADY,
          AXI_STR_TXD_TLAST      => AXI_STR_TXD_TLAST,
          AXI_STR_TXD_TSTRB      => AXI_STR_TXD_TSTRB,
          AXI_STR_TXD_TDATA      => AXI_STR_TXD_TDATA,
          -- AXI Stream Control signals
          AXI_STR_TXC_ACLK       => AXI_STR_TXC_ACLK,
          reset2axi_str_txc      => reset2axi_str_txc,
          AXI_STR_TXC_TVALID     => AXI_STR_TXC_TVALID,
          AXI_STR_TXC_TREADY     => AXI_STR_TXC_TREADY,
          AXI_STR_TXC_TLAST      => AXI_STR_TXC_TLAST,
          AXI_STR_TXC_TSTRB      => AXI_STR_TXC_TSTRB,
          AXI_STR_TXC_TDATA      => AXI_STR_TXC_TDATA,

          -- Write Port - AXI Stream TxData
          Axi_Str_TxD_2_Mem_Din  => Axi_Str_TxD_2_Mem_Din,       --: out std_logic_vector(c_TxD_write_width_b-1 downto 0);
          Axi_Str_TxD_2_Mem_Addr => Axi_Str_TxD_2_Mem_Addr,      --: out std_logic_vector(c_TxD_addrb_width-1   downto 0);
          Axi_Str_TxD_2_Mem_En   => Axi_Str_TxD_2_Mem_En,        --: out std_logic := '1';
          Axi_Str_TxD_2_Mem_We   => Axi_Str_TxD_2_Mem_We,        --: out std_logic_vector(c_TxD_web_width-1     downto 0);
          Axi_Str_TxD_2_Mem_Dout => Axi_Str_TxD_2_Mem_Dout,      --: in  std_logic_vector(c_TxD_read_width_b-1  downto 0);

          -- Write Port - AXI Stream TxControl
          Axi_Str_TxC_2_Mem_Din  => Axi_Str_TxC_2_Mem_Din,       --: out std_logic_vector(c_TxD_write_width_b-1 downto 0);
          Axi_Str_TxC_2_Mem_Addr => Axi_Str_TxC_2_Mem_Addr,      --: out std_logic_vector(c_TxD_addrb_width-1   downto 0);
          Axi_Str_TxC_2_Mem_En   => Axi_Str_TxC_2_Mem_En,        --: out std_logic := '1';
          Axi_Str_TxC_2_Mem_We   => Axi_Str_TxC_2_Mem_We,        --: out std_logic_vector(c_TxD_web_width-1     downto 0);
          Axi_Str_TxC_2_Mem_Dout => Axi_Str_TxC_2_Mem_Dout,      --: in  std_logic_vector(c_TxD_read_width_b-1  downto 0);

          tx_vlan_bram_addr      => tx_vlan_bram_addr,
          tx_vlan_bram_din       => tx_vlan_bram_din,
          tx_vlan_bram_en        => tx_vlan_bram_en,

          enable_newFncEn        => enable_newFncEn,
          transMode_cross        => transMode_cross,
          tagMode_cross          => tagMode_cross,
          strpMode_cross         => strpMode_cross,

          tpid0_cross            => tpid0_cross,
          tpid1_cross            => tpid1_cross,
          tpid2_cross            => tpid2_cross,
          tpid3_cross            => tpid3_cross,

          newTagData_cross       => newTagData_cross,

          tx_init_in_prog        => tx_init_in_prog

        );


       TX_MEM_INTERFACE : tx_mem_if
       --BRAM between AXI Stream Interface and Tx Client Interface
       generic map(
          C_FAMILY                 => C_FAMILY,

          -- Read Port - AXI Stream TxData
          c_TxD_write_width_a      => c_TxD_write_width_a,
          c_TxD_read_width_a       => c_TxD_read_width_a,
          c_TxD_write_depth_a      => c_TxD_write_depth_a,
          c_TxD_read_depth_a       => c_TxD_read_depth_a,
          c_TxD_addra_width        => c_TxD_addra_width,
          c_TxD_wea_width          => c_TxD_wea_width,
          -- Write Port - AXI Stream TxData
          c_TxD_write_width_b      => c_TxD_write_width_b,
          c_TxD_read_width_b       => c_TxD_read_width_b,
          c_TxD_write_depth_b      => c_TxD_write_depth_b,
          c_TxD_read_depth_b       => c_TxD_read_depth_b,
          c_TxD_addrb_width        => c_TxD_addrb_width,
          c_TxD_web_width          => c_TxD_web_width,

          -- Read Port - AXI Stream TxControl
          c_TxC_write_width_a      => c_TxC_write_width_a,
          c_TxC_read_width_a       => c_TxC_read_width_a,
          c_TxC_write_depth_a      => c_TxC_write_depth_a,
          c_TxC_read_depth_a       => c_TxC_read_depth_a,
          c_TxC_addra_width        => c_TxC_addra_width,
          c_TxC_wea_width          => c_TxC_wea_width,
          -- Write Port - AXI Stream TxControl
          c_TxC_write_width_b      => c_TxC_write_width_b,
          c_TxC_read_width_b       => c_TxC_read_width_b,
          c_TxC_write_depth_b      => c_TxC_write_depth_b,
          c_TxC_read_depth_b       => c_TxC_read_depth_b,
          c_TxC_addrb_width        => c_TxC_addrb_width,
          c_TxC_web_width          => c_TxC_web_width

        )
        port map  (
          -- Read Port - AXI Stream TxData
          TX_CLIENT_CLK             => tx_mac_aclk,            --: in  std_logic;
          reset2tx_client           => tx_reset,          --: in  std_logic;
          Tx_Client_TxD_2_Mem_Din   => Tx_Client_TxD_2_Mem_Din,  --: in  std_logic_vector(c_TxD_write_width_a-1 downto 0);
          Tx_Client_TxD_2_Mem_Addr  => Tx_Client_TxD_2_Mem_Addr, --: in  std_logic_vector(c_TxD_addra_width-1   downto 0);
          Tx_Client_TxD_2_Mem_En    => Tx_Client_TxD_2_Mem_En,   --: in  std_logic := '1';
          Tx_Client_TxD_2_Mem_We    => Tx_Client_TxD_2_Mem_We,   --: in  std_logic_vector(c_TxD_wea_width-1     downto 0);
          Tx_Client_TxD_2_Mem_Dout  => Tx_Client_TxD_2_Mem_Dout, --: out std_logic_vector(c_TxD_read_width_a-1  downto 0);
          -- Write Port - AXI Stream TxData
          AXI_STR_TXD_ACLK          => AXI_STR_TXD_ACLK,         --: in  std_logic := '0';
          reset2axi_str_txd         => reset2axi_str_txd,        --: in  std_logic;
          Axi_Str_TxD_2_Mem_Din     => Axi_Str_TxD_2_Mem_Din,    --: in  std_logic_vector(c_TxD_write_width_b-1 downto 0);
          Axi_Str_TxD_2_Mem_Addr    => Axi_Str_TxD_2_Mem_Addr,   --: in  std_logic_vector(c_TxD_addrb_width-1   downto 0);
          Axi_Str_TxD_2_Mem_En      => Axi_Str_TxD_2_Mem_En,     --: in  std_logic := '1';
          Axi_Str_TxD_2_Mem_We      => Axi_Str_TxD_2_Mem_We,     --: in  std_logic_vector(c_TxD_web_width-1     downto 0);
          Axi_Str_TxD_2_Mem_Dout    => Axi_Str_TxD_2_Mem_Dout,   --: out std_logic_vector(c_TxD_read_width_b-1  downto 0);

          -- Read Port - AXI Stream TxControl
          Tx_Client_TxC_2_Mem_Din   => Tx_Client_TxC_2_Mem_Din,  --: in  std_logic_vector(c_TxD_write_width_a-1 downto 0);
          Tx_Client_TxC_2_Mem_Addr  => Tx_Client_TxC_2_Mem_Addr, --: in  std_logic_vector(c_TxD_addra_width-1   downto 0);
          Tx_Client_TxC_2_Mem_En    => Tx_Client_TxC_2_Mem_En,   --: in  std_logic := '1';
          Tx_Client_TxC_2_Mem_We    => Tx_Client_TxC_2_Mem_We,   --: in  std_logic_vector(c_TxD_wea_width-1     downto 0);
          Tx_Client_TxC_2_Mem_Dout  => Tx_Client_TxC_2_Mem_Dout, --: out std_logic_vector(c_TxD_read_width_a-1  downto 0);
          -- Write Port - AXI Stream TxControl
          AXI_STR_TXC_ACLK          => AXI_STR_TXC_ACLK,         --: in  std_logic := '0';
          reset2axi_str_txc         => reset2axi_str_txc,        --: in  std_logic;
          Axi_Str_TxC_2_Mem_Din     => Axi_Str_TxC_2_Mem_Din,    --: in  std_logic_vector(c_TxD_write_width_b-1 downto 0);
          Axi_Str_TxC_2_Mem_Addr    => Axi_Str_TxC_2_Mem_Addr,   --: in  std_logic_vector(c_TxD_addrb_width-1   downto 0);
          Axi_Str_TxC_2_Mem_En      => Axi_Str_TxC_2_Mem_En,     --: in  std_logic := '1';
          Axi_Str_TxC_2_Mem_We      => Axi_Str_TxC_2_Mem_We,     --: in  std_logic_vector(c_TxD_web_width-1     downto 0);
          Axi_Str_TxC_2_Mem_Dout    => Axi_Str_TxC_2_Mem_Dout    --: out std_logic_vector(c_TxD_read_width_b-1  downto 0);
        );

GEN_1G_MAC_IF: if (C_SPEED_2P5 = 0) generate 
begin
        TX_EMAC_INTERFACE : tx_emac_if
        --  Interface for Transmit AxiStream Data and Control; and Tx Memory
        generic map (
          C_FAMILY                  => C_FAMILY,                 --: string                        := "virtex6";
          C_HALFDUP                 => C_HALFDUP,                --: integer range 0 to 1          := 0;
          C_TXMEM                   => C_TXMEM,                  --: integer                       := 4096;
          C_TXCSUM                  => C_TXCSUM,                 --: integer range 0 to 2          := 0;
          C_ENABLE_1588             => C_ENABLE_1588,

          -- Read Port - AXI Stream TxData
          c_TxD_write_width_a       => c_TxD_write_width_a,
          c_TxD_read_width_a        => c_TxD_read_width_a,
          c_TxD_write_depth_a       => c_TxD_write_depth_a,
          c_TxD_read_depth_a        => c_TxD_read_depth_a,
          c_TxD_addra_width         => c_TxD_addra_width,
          c_TxD_wea_width           => c_TxD_wea_width,

          -- Read Port - AXI Stream TxControl
          c_TxC_write_width_a       => c_TxC_write_width_a,
          c_TxC_read_width_a        => c_TxC_read_width_a,
          c_TxC_write_depth_a       => c_TxC_write_depth_a,
          c_TxC_read_depth_a        => c_TxC_read_depth_a,
          c_TxC_addra_width         => c_TxC_addra_width,
          c_TxC_wea_width           => c_TxC_wea_width,

          c_TxD_addrb_width         => c_TxD_addrb_width
        )
        port map  (
          tx_client_10_100          => tx_client_10_100,

          -- Read Port - AXI Stream TxData
          reset2tx_client           => tx_reset,          --: in  std_logic;
          Tx_Client_TxD_2_Mem_Din   => Tx_Client_TxD_2_Mem_Din,  --: out std_logic_vector(c_TxD_write_width_a-1 downto 0);
          Tx_Client_TxD_2_Mem_Addr  => Tx_Client_TxD_2_Mem_Addr, --: out std_logic_vector(c_TxD_addra_width-1   downto 0);
          Tx_Client_TxD_2_Mem_En    => Tx_Client_TxD_2_Mem_En,   --: out std_logic := '1';
          Tx_Client_TxD_2_Mem_We    => Tx_Client_TxD_2_Mem_We,   --: out std_logic_vector(c_TxD_wea_width-1     downto 0);
          Tx_Client_TxD_2_Mem_Dout  => Tx_Client_TxD_2_Mem_Dout, --: in  std_logic_vector(c_TxD_read_width_a-1  downto 0);

          -- Read Port - AXI Stream TxControl
          reset2axi_str_txd         => reset2axi_str_txd,        --: in  std_logic;
          Tx_Client_TxC_2_Mem_Din   => Tx_Client_TxC_2_Mem_Din,  --: out std_logic_vector(c_TxD_write_width_a-1 downto 0);
          Tx_Client_TxC_2_Mem_Addr  => Tx_Client_TxC_2_Mem_Addr, --: out std_logic_vector(c_TxD_addra_width-1   downto 0);
          Tx_Client_TxC_2_Mem_En    => Tx_Client_TxC_2_Mem_En,   --: out std_logic := '1';
          Tx_Client_TxC_2_Mem_We    => Tx_Client_TxC_2_Mem_We,   --: out std_logic_vector(c_TxD_wea_width-1     downto 0);
          Tx_Client_TxC_2_Mem_Dout  => Tx_Client_TxC_2_Mem_Dout, --: in  std_logic_vector(c_TxD_read_width_a-1  downto 0);


          tx_axi_clk                => tx_mac_aclk,
          tx_reset_out              => tx_reset,
          tx_axis_mac_tdata         => tx_axis_mac_tdata_int , --tx_axis_mac_tdata,
          tx_axis_mac_tvalid        => tx_axis_mac_tvalid_int, --tx_axis_mac_tvalid,
          tx_axis_mac_tlast         => tx_axis_mac_tlast_int , --tx_axis_mac_tlast,
          tx_axis_mac_tuser         => tx_axis_mac_tuser_int , --tx_axis_mac_tuser,
          tx_axis_mac_tready        => tx_axis_mac_tready_int, --tx_axis_mac_tready,
          tx_collision              => tx_collision,           --tx_collision,
          tx_retransmit             => tx_retransmit,          --tx_retransmit,

          tx_cmplt                  => tx_cmplt,

          tx_init_in_prog_cross     => tx_init_in_prog_cross
        );

end generate GEN_1G_MAC_IF;

GEN_2P5G_MAC_IF: if (C_SPEED_2P5 = 1) generate 
begin
        TX_EMAC_INTERFACE : tx_emac_if_2g5
        --  Interface for Transmit AxiStream Data and Control; and Tx Memory
        generic map (
          C_FAMILY                  => C_FAMILY,                 --: string                        := "virtex6";
          C_HALFDUP                 => C_HALFDUP,                --: integer range 0 to 1          := 0;
          C_TXMEM                   => C_TXMEM,                  --: integer                       := 4096;
          C_TXCSUM                  => C_TXCSUM,                 --: integer range 0 to 2          := 0;
          C_ENABLE_1588             => C_ENABLE_1588,

          -- Read Port - AXI Stream TxData
          c_TxD_write_width_a       => c_TxD_write_width_a,
          c_TxD_read_width_a        => c_TxD_read_width_a,
          c_TxD_write_depth_a       => c_TxD_write_depth_a,
          c_TxD_read_depth_a        => c_TxD_read_depth_a,
          c_TxD_addra_width         => c_TxD_addra_width,
          c_TxD_wea_width           => c_TxD_wea_width,

          -- Read Port - AXI Stream TxControl
          c_TxC_write_width_a       => c_TxC_write_width_a,
          c_TxC_read_width_a        => c_TxC_read_width_a,
          c_TxC_write_depth_a       => c_TxC_write_depth_a,
          c_TxC_read_depth_a        => c_TxC_read_depth_a,
          c_TxC_addra_width         => c_TxC_addra_width,
          c_TxC_wea_width           => c_TxC_wea_width,

          c_TxD_addrb_width         => c_TxD_addrb_width
        )
        port map  (
          tx_client_10_100          => tx_client_10_100,

          -- Read Port - AXI Stream TxData
          reset2tx_client           => tx_reset,          --: in  std_logic;
          Tx_Client_TxD_2_Mem_Din   => Tx_Client_TxD_2_Mem_Din,  --: out std_logic_vector(c_TxD_write_width_a-1 downto 0);
          Tx_Client_TxD_2_Mem_Addr  => Tx_Client_TxD_2_Mem_Addr, --: out std_logic_vector(c_TxD_addra_width-1   downto 0);
          Tx_Client_TxD_2_Mem_En    => Tx_Client_TxD_2_Mem_En,   --: out std_logic := '1';
          Tx_Client_TxD_2_Mem_We    => Tx_Client_TxD_2_Mem_We,   --: out std_logic_vector(c_TxD_wea_width-1     downto 0);
          Tx_Client_TxD_2_Mem_Dout  => Tx_Client_TxD_2_Mem_Dout, --: in  std_logic_vector(c_TxD_read_width_a-1  downto 0);

          -- Read Port - AXI Stream TxControl
          reset2axi_str_txd         => reset2axi_str_txd,        --: in  std_logic;
          Tx_Client_TxC_2_Mem_Din   => Tx_Client_TxC_2_Mem_Din,  --: out std_logic_vector(c_TxD_write_width_a-1 downto 0);
          Tx_Client_TxC_2_Mem_Addr  => Tx_Client_TxC_2_Mem_Addr, --: out std_logic_vector(c_TxD_addra_width-1   downto 0);
          Tx_Client_TxC_2_Mem_En    => Tx_Client_TxC_2_Mem_En,   --: out std_logic := '1';
          Tx_Client_TxC_2_Mem_We    => Tx_Client_TxC_2_Mem_We,   --: out std_logic_vector(c_TxD_wea_width-1     downto 0);
          Tx_Client_TxC_2_Mem_Dout  => Tx_Client_TxC_2_Mem_Dout, --: in  std_logic_vector(c_TxD_read_width_a-1  downto 0);


          tx_axi_clk                => tx_mac_aclk,
          tx_reset_out              => tx_reset,
          tx_axis_mac_tdata         => tx_axis_mac_tdata_int , --tx_axis_mac_tdata,
          tx_axis_mac_tvalid        => tx_axis_mac_tvalid_int, --tx_axis_mac_tvalid,
          tx_axis_mac_tlast         => tx_axis_mac_tlast_int , --tx_axis_mac_tlast,
          tx_axis_mac_tuser         => tx_axis_mac_tuser_int , --tx_axis_mac_tuser,
          tx_axis_mac_tready        => tx_axis_mac_tready_int, --tx_axis_mac_tready,
          tx_collision              => tx_collision,           --tx_collision,
          tx_retransmit             => tx_retransmit,          --tx_retransmit,

          tx_cmplt                  => tx_cmplt,

          tx_init_in_prog_cross     => tx_init_in_prog_cross
        );
          
end generate GEN_2P5G_MAC_IF;
          tx_axis_mac_tvalid     <= tx_axis_mac_tvalid_int;
          tx_axis_mac_tlast      <= tx_axis_mac_tlast_int;
          tx_axis_mac_tuser      <= tx_axis_mac_tuser_int;
          tx_axis_mac_tready_int <= tx_axis_mac_tready;
          tx_axis_mac_tdata      <= tx_axis_mac_tdata_int;

end imp;


------------------------------------------------------------------------------
-- registers - entity and arch
------------------------------------------------------------------------------
--
-- DISCLAIMER OF LIABILITY
--
-- This file contains proprietary and confidential information of

-- from Xilinx, and may be used, copied and/or disclosed only

--
-- XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
-- ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
-- EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
-- LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
-- MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
-- does not warrant that functions included in the Materials will

-- Materials will be uninterrupted or error-free, or that defects
-- in the Materials will be corrected. Furthermore, Xilinx does
-- not warrant or make any representations regarding use, or the
-- results of the use, of the Materials in terms of correctness,
-- accuracy, reliability or otherwise.
--
-- Xilinx products are not designed or intended to be fail-safe,
-- or for use in any application requiring fail-safe performance,
-- such as life-support or safety devices or systems, Class III
-- medical devices, nuclear facilities, applications related to
-- the deployment of airbags, or any other applications that could
-- lead to death, personal injury or severe property or
-- environmental damage (individually and collectively, "critical
-- applications"). Customer assumes the sole risk and liability
-- of any use of Xilinx products in critical applications,
-- subject only to applicable laws and regulations governing
-- limitations on product liability.
--
-- Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
-- All rights reserved.
--
-- This disclaimer and copyright notice must be retained as part
-- of this file at all times.
--

------------------------------------------------------------------------------
-- Filename:        registers.vhd
-- Version:         v2.00a
-- Description:     Include a meaningful description of your file. Multi-line
--                  descriptions should align with each other
--
--  Addr   REG    Chipselect #
-- offset
-- 0x000   RAF   Bus2IP_Wr/RdCE(0) Bus2IP_CS(0)
-- 0x004   TPF   Bus2IP_Wr/RdCE(1) Bus2IP_CS(0)
-- 0x008   IFGP  Bus2IP_Wr/RdCE(2) Bus2IP_CS(0)
-- 0x00C   IS    Bus2IP_Wr/RdCE(3) Bus2IP_CS(0)
-- 0x010   IP    Bus2IP_Wr/RdCE(4) Bus2IP_CS(0)
-- 0x014   IE    Bus2IP_Wr/RdCE(5) Bus2IP_CS(0)
-- 0x018   TTAG  Bus2IP_Wr/RdCE(6) Bus2IP_CS(0)
-- 0x01C   RTAG  Bus2IP_Wr/RdCE(7) Bus2IP_CS(0)
-- 0x020   UAWL  Bus2IP_Wr/RdCE(8)  Bus2IP_CS(0)
-- 0x024   UAWU  Bus2IP_Wr/RdCE(9)  Bus2IP_CS(0)
-- 0x028   TPID0 Bus2IP_Wr/RdCE(10) Bus2IP_CS(0)
-- 0x02C   TPID1 Bus2IP_Wr/RdCE(11) Bus2IP_CS(0)
--
-- 0x0000200 - 0x00007FC stats & temac regs  Bus2IP_Wr/RdCE(16) Bus2IP_CS(1)
-- 0x0004000 - 0x0007FFC TX VLAN TRANS  BRAM Bus2IP_Wr/RdCE(17) Bus2IP_CS(2)
-- 0x0008000 - 0x000BFFC RX VLAN TRANS  BRAM Bus2IP_Wr/RdCE(18) Bus2IP_CS(3)
-- 0x0010000 - 0x0013FFC AVB                 Bus2IP_Wr/RdCE(19) Bus2IP_CS(4)
-- 0x0020000 - 0x003FFFC Multicast ADDR BRAM Bus2IP_Wr/RdCE(20) Bus2IP_CS(5)
--
------------------------------------------------------------------------------
-- Structure:   This section should show the hierarchical structure of the
--              designs. Separate lines with blank lines if necessary to improve
--              readability.
--
--              top_level.vhd
--                  -- second_level_file1.vhd
--                      -- third_level_file1.vhd
--                          -- fourth_level_file.vhd
--                      -- third_level_file2.vhd
--                  -- second_level_file2.vhd
--                  -- second_level_file3.vhd
--
--              This section is optional for common/shared modules but should
--              contain a statement stating it is a common/shared module.
------------------------------------------------------------------------------
-- Author:
-- History:
--
--
------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      AxiReset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_cmb"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.registers_pack.all;

--library lib_bmg_v1_0;
--use lib_bmg_v1_0.all;

Library xpm;
use xpm.vcomponents.all;

entity registers is
  generic
  (
    C_FAMILY       : string   := "virtex5";
    C_TXVLAN_TRAN  : integer  := 1;
    C_TXVLAN_TAG   : integer  := 1;
    C_TXVLAN_STRP  : integer  := 1;
    C_RXVLAN_TRAN  : integer  := 1;
    C_RXVLAN_TAG   : integer  := 1;
    C_RXVLAN_STRP  : integer  := 1;
    C_MCAST_EXTEND : integer  := 1;
    C_TXVLAN_WIDTH : integer  := 1;
    C_RXVLAN_WIDTH : integer  := 1
  );
  port
  (
    AxiClk                    : in  std_logic;                    --  AXI4-Lite Clock
    AXI_STR_TXD_ACLK          : in  std_logic;                    --  AXI-Stream Transmit Data Clock
    RxClClk                   : in  std_logic;                    --  Receive Client Clock
    AxiReset                  : in  std_logic;                    --  AXI4-Lite Reset
    IP2Bus_Data               : out std_logic_vector(0 to 31);    --  AXI Ethernet to AXI4-Lite Data
    IP2Bus_WrAck              : out std_logic;                    --  AXI Ethernet to AXI4-Lite Write Ack
    IP2Bus_RdAck              : out std_logic;                    --  AXI Ethernet to AXI4-Lite Read Ack
    Bus2IP_Addr               : in  std_logic_vector(0 to 31);    --  AXI4-Lite to AXI Ethernet Addr
    Bus2IP_Data               : in  std_logic_vector(0 to 31);    --  AXI4-Lite to AXI Ethernet Data
    Bus2IP_RNW                : in  std_logic;                    --  AXI4-Lite to AXI Ethernet RNW
    Bus2IP_CS                 : in  std_logic_vector(0 to 10);    --  AXI4-Lite to AXI Ethernet CS
    Bus2IP_RdCE               : in  std_logic_vector(0 to 41);    --  AXI4-Lite to AXI Ethernet RdCE
    Bus2IP_WrCE               : in  std_logic_vector(0 to 41);    --  AXI4-Lite to AXI Ethernet WrCE
    IntrptsIn                 : in  std_logic_vector(23 to 31);   --  Interrupts in
    TPReq                     : out std_logic;                    --  Transmit Pause Request
    CrRegData                 : out std_logic_vector(17 to 31);   --  RAF Register
    TpRegData                 : out std_logic_vector(16 to 31);   --  Transmit Pause Data
    IfgpRegData               : out std_logic_vector(24 to 31);   --  Inter Frame Gap Data
    IsRegData                 : out std_logic_vector(23 to 31);   --  Interrupt Status Register
    IpRegData                 : out std_logic_vector(23 to 31);   --  Interrupt Pending Register
    IeRegData                 : out std_logic_vector(23 to 31);   --  Interrupt Enable Register
    IntrptOut                 : out std_logic;                    --  Interrupt Out
    TtagRegData               : out std_logic_vector(0 to 31);    --  Transmit Tag Register
    RtagRegData               : out std_logic_vector(0 to 31);    --  Receive Tag Register
    Tpid0RegData              : out std_logic_vector(0 to 31);    --  VLAN TPID Reg 0
    Tpid1RegData              : out std_logic_vector(0 to 31);    --  VLAN TPID Reg 1
    pcspma_status_cross       : in  std_logic_vector(16 to 31);   --  PCS PMA Link Status Vector
    UawLRegData               : out std_logic_vector(0 to 31);    --  Unicast Address Word Lower
    UawURegData               : out std_logic_vector(16 to 31);   --  Unicast Address Word Upper
    RxClClkMcastAddr          : in  std_logic_vector(0 to 14);    --  Receive Extended Multicast Address
    RxClClkMcastEn            : in  std_logic;                    --  Receive Extended Multicast Enable
    RxClClkMcastRdData        : out std_logic_vector(0 to 0);     --  Receive Extended Multicast Data
    AxiStrTxDClkTxVlanAddr    : in  std_logic_vector(0 to 11);    --  Transmit VLAN BRAM Addr
    AxiStrTxDClkTxVlanRdData  : out std_logic_vector(18 to 31);   --  Transmit VLAN BRAM Read Data
    RxClClkRxVlanAddr         : in  std_logic_vector(0 to 11);    --  Receive VLAN BRAM Addr
    RxClClkRXVlanRdData       : out std_logic_vector(18 to 31);   --  Receive VLAN BRAM Read Data
    AxiStrTxDClkTxVlanBramEnA : in  std_logic;                    --  Transmit VLAN BRAM Enable
    RxClClkRxVlanBramEnA      : in  std_logic                     --  Receive VLAN BRAM Enable
  );
end registers;

architecture imp of registers is

signal crRdData      : std_logic_vector(17 to 31);
signal tpRdData      : std_logic_vector(16 to 31);
signal ifgpRdData    : std_logic_vector(24 to 31);
signal isRdData      : std_logic_vector(23 to 31);
signal ieRdData      : std_logic_vector(23 to 31);
signal ipRdData      : std_logic_vector(23 to 31);
signal ttagRdData    : std_logic_vector(0 to 31);
signal rtagRdData    : std_logic_vector(0 to 31);
signal tpid0RdData   : std_logic_vector(0 to 31);
signal tpid1RdData   : std_logic_vector(0 to 31);
signal pcspma_status : std_logic_vector(16 to 31);
signal uawLRdData    : std_logic_vector(0 to 31);
signal uawURdData    : std_logic_vector(16 to 31);

signal isRegData_i   : std_logic_vector(23 to 31);
signal ieRegData_i   : std_logic_vector(23 to 31);
signal ttagRegData_i : std_logic_vector(0 to 31);
signal rtagRegData_i : std_logic_vector(0 to 31);
signal tpid0RegData_i: std_logic_vector(0 to 31);
signal tpid1RegData_i: std_logic_vector(0 to 31);
signal uawLRegData_i : std_logic_vector(0 to 31);
signal uawURegData_i : std_logic_vector(16 to 31);
signal axiClkMcastRdData    : std_logic_vector(0 to 0);
signal axiClkMcastRdData_i  : std_logic_vector(0 to 0);
signal axiClkTxVlanRdData   : std_logic_vector(18 to 31);
signal axiClkTxVlanRdData_i : std_logic_vector(((31-C_TXVLAN_WIDTH)+1) to 31);
signal axiClkTxVlanWrData_i : std_logic_vector(((31-C_TXVLAN_WIDTH)+1) to 31);
signal axiClkRxVlanRdData   : std_logic_vector(18 to 31);
signal axiClkRxVlanRdData_i : std_logic_vector(((31-C_RXVLAN_WIDTH)+1) to 31);
signal axiClkRxVlanWrData_i : std_logic_vector(((31-C_RXVLAN_WIDTH)+1) to 31);
signal AxiStrTxDClkTxRdData_i   : std_logic_vector(((31-C_TXVLAN_WIDTH)+1) to 31);
signal rxClClkRxRdData_i   : std_logic_vector(((31-C_RXVLAN_WIDTH)+1) to 31);
signal txvlan_dina    : std_logic_vector(((31-C_TXVLAN_WIDTH)+1) to 31);
signal rxvlan_dina    : std_logic_vector(((31-C_RXVLAN_WIDTH)+1) to 31);
signal rdData          : std_logic_vector(0 to 31);
signal softRead        : std_logic;
signal softWrite       : std_logic;
signal temacDcr_DBus_i : std_logic_vector(0 to 31);
signal softRead_d1     : std_logic;
signal softWrite_d1    : std_logic;

signal iP2Bus_WrAck_i  : std_logic;
signal iP2Bus_RdAck_i  : std_logic;

signal rdAckBlocker    : std_logic;
signal wrAckBlocker    : std_logic;

signal bus2IP_WrCE_17_d1 : std_logic;
signal bus2IP_WrCE_17_en : std_logic;

signal bus2IP_WrCE_18_d1 : std_logic;
signal bus2IP_WrCE_18_en : std_logic;

signal bus2IP_WrCE_20_d1 : std_logic;
signal bus2IP_WrCE_20_en : std_logic;

signal zeroes            : std_logic_vector(23 downto 0);

begin
  PIPE_RAM_WRITE_PROCESS: process (AxiClk)
  begin
    if (AxiClk'event and AxiClk = '1') then
      if (AxiReset = '1') then
        bus2IP_WrCE_17_d1     <= '0';
        bus2IP_WrCE_17_en     <= '0';
        bus2IP_WrCE_18_d1     <= '0';
        bus2IP_WrCE_18_en     <= '0';
        bus2IP_WrCE_20_d1     <= '0';
        bus2IP_WrCE_20_en     <= '0';
      else
        bus2IP_WrCE_17_d1     <= Bus2IP_WrCE(17);
        bus2IP_WrCE_17_en     <= Bus2IP_WrCE(17) and not(bus2IP_WrCE_17_d1);
        bus2IP_WrCE_18_d1     <= Bus2IP_WrCE(18);
        bus2IP_WrCE_18_en     <= Bus2IP_WrCE(18) and not(bus2IP_WrCE_18_d1);
        bus2IP_WrCE_20_d1     <= Bus2IP_WrCE(20);
        bus2IP_WrCE_20_en     <= Bus2IP_WrCE(20) and not(bus2IP_WrCE_20_d1);
      end if;
    end if;
  end process;

  txvlan_dina <= (others => '0');
  rxvlan_dina <= (others => '0');

  -- TX VLAN --
  TX_VLAN_TRAN_STRP_TAG : if (C_TXVLAN_TRAN = 1 and C_TXVLAN_STRP = 1 and C_TXVLAN_TAG = 1) generate
  begin
    axiClkTxVlanRdData   <= axiClkTxVlanRdData_i when (Bus2IP_RdCE(17) = '1') else (others => '0');
    axiClkTxVlanWrData_i <= Bus2IP_Data(18 to 31);
    AxiStrTxDClkTxVlanRdData  <= AxiStrTxDClkTxRdData_i;
  end generate TX_VLAN_TRAN_STRP_TAG;

  TX_VLAN_TRAN_STRP : if (C_TXVLAN_TRAN = 1 and C_TXVLAN_STRP = 1 and C_TXVLAN_TAG = 0) generate
  begin
    axiClkTxVlanRdData   <= axiClkTxVlanRdData_i & '0' when (Bus2IP_RdCE(17) = '1') else (others => '0');
    axiClkTxVlanWrData_i <= Bus2IP_Data(18 to 30);
    AxiStrTxDClkTxVlanRdData  <= AxiStrTxDClkTxRdData_i & '0';
  end generate TX_VLAN_TRAN_STRP;

  TX_VLAN_TRAN_TAG : if (C_TXVLAN_TRAN = 1 and C_TXVLAN_STRP = 0 and C_TXVLAN_TAG = 1) generate
  begin
    axiClkTxVlanRdData   <= axiClkTxVlanRdData_i(19 to 30) & '0' & axiClkTxVlanRdData_i(31)
                              when (Bus2IP_RdCE(17) = '1') else (others => '0');
    axiClkTxVlanWrData_i <= Bus2IP_Data(18 to 29)& Bus2IP_Data(31);
    AxiStrTxDClkTxVlanRdData  <= AxiStrTxDClkTxRdData_i(19 to 30) & '0' & AxiStrTxDClkTxRdData_i(31);
  end generate TX_VLAN_TRAN_TAG;

  TX_VLAN_TRAN : if (C_TXVLAN_TRAN = 1 and C_TXVLAN_STRP = 0 and C_TXVLAN_TAG = 0) generate
  begin
    axiClkTxVlanRdData   <= axiClkTxVlanRdData_i(20 to 31) & "00" when (Bus2IP_RdCE(17) = '1') else (others => '0');
    axiClkTxVlanWrData_i <= Bus2IP_Data(18 to 29);
    AxiStrTxDClkTxVlanRdData  <= AxiStrTxDClkTxRdData_i(20 to 31) & "00";
  end generate TX_VLAN_TRAN;

  TX_VLAN_STRP_TAG : if (C_TXVLAN_TRAN = 0 and C_TXVLAN_STRP = 1 and C_TXVLAN_TAG = 1) generate
  begin
    axiClkTxVlanRdData   <= "000000000000" & axiClkTxVlanRdData_i when (Bus2IP_RdCE(17) = '1') else (others => '0');
    axiClkTxVlanWrData_i <= Bus2IP_Data(30 to 31);
    AxiStrTxDClkTxVlanRdData  <= "000000000000" & AxiStrTxDClkTxRdData_i;
  end generate TX_VLAN_STRP_TAG;

  TX_VLAN_STRP : if (C_TXVLAN_TRAN = 0 and C_TXVLAN_STRP = 1 and C_TXVLAN_TAG = 0) generate
  begin
    axiClkTxVlanRdData   <= "000000000000" & axiClkTxVlanRdData_i & '0'
                              when (Bus2IP_RdCE(17) = '1') else (others => '0');
    axiClkTxVlanWrData_i <= Bus2IP_Data(30 to 30);
    AxiStrTxDClkTxVlanRdData  <= "000000000000" & AxiStrTxDClkTxRdData_i & '0';
  end generate TX_VLAN_STRP;

  TX_VLAN_TAG : if (C_TXVLAN_TRAN = 0 and C_TXVLAN_STRP = 0 and C_TXVLAN_TAG = 1) generate
  begin
    axiClkTxVlanRdData   <= "000000000000" & '0' & axiClkTxVlanRdData_i
                              when (Bus2IP_RdCE(17) = '1') else (others => '0');
    axiClkTxVlanWrData_i <= Bus2IP_Data(31 to 31);
    AxiStrTxDClkTxVlanRdData  <= "000000000000" & '0' & AxiStrTxDClkTxRdData_i;
  end generate TX_VLAN_TAG;

  TX_VLAN_NONE : if (C_TXVLAN_TRAN = 0 and C_TXVLAN_STRP = 0 and C_TXVLAN_TAG = 0) generate
  begin
    axiClkTxVlanRdData   <= (others => '0');
    AxiStrTxDClkTxVlanRdData  <= (others => '0');
  end generate TX_VLAN_NONE;

  -- RX VLAN --
  RX_VLAN_TRAN_STRP_TAG : if (C_RXVLAN_TRAN = 1 and C_RXVLAN_STRP = 1 and C_RXVLAN_TAG = 1) generate
  begin
    axiClkRXVlanRdData    <= axiClkRXVlanRdData_i when (Bus2IP_RdCE(18) = '1') else (others => '0');
    axiClkRXVlanWrData_i  <= Bus2IP_Data(18 to 31);
    RxClClkRXVlanRdData   <= rxClClkRxRdData_i;
  end generate RX_VLAN_TRAN_STRP_TAG;

  RX_VLAN_TRAN_STRP : if (C_RXVLAN_TRAN = 1 and C_RXVLAN_STRP = 1 and C_RXVLAN_TAG = 0) generate
  begin
    axiClkRXVlanRdData    <= axiClkRXVlanRdData_i & '0' when (Bus2IP_RdCE(18) = '1') else (others => '0');
    axiClkRXVlanWrData_i  <= Bus2IP_Data(18 to 30);
    RxClClkRXVlanRdData   <= rxClClkRxRdData_i & '0';
  end generate RX_VLAN_TRAN_STRP;

  RX_VLAN_TRAN_TAG : if (C_RXVLAN_TRAN = 1 and C_RXVLAN_STRP = 0 and C_RXVLAN_TAG = 1) generate
  begin
    axiClkRXVlanRdData    <= axiClkRXVlanRdData_i(19 to 30) & '0' & axiClkRXVlanRdData_i(31)
                              when (Bus2IP_RdCE(18) = '1') else (others => '0');
    axiClkRXVlanWrData_i  <= Bus2IP_Data(18 to 29)& Bus2IP_Data(31);
    RxClClkRXVlanRdData   <= rxClClkRxRdData_i(19 to 30) & '0' & rxClClkRxRdData_i(31);
  end generate RX_VLAN_TRAN_TAG;

  RX_VLAN_TRAN : if (C_RXVLAN_TRAN = 1 and C_RXVLAN_STRP = 0 and C_RXVLAN_TAG = 0) generate
  begin
    axiClkRXVlanRdData    <= axiClkRXVlanRdData_i(20 to 31) & "00" when (Bus2IP_RdCE(18) = '1') else (others => '0');
    axiClkRXVlanWrData_i  <= Bus2IP_Data(18 to 29);
    RxClClkRXVlanRdData   <= rxClClkRxRdData_i(20 to 31) & "00";
  end generate RX_VLAN_TRAN;

  RX_VLAN_STRP_TAG : if (C_RXVLAN_TRAN = 0 and C_RXVLAN_STRP = 1 and C_RXVLAN_TAG = 1) generate
  begin
    axiClkRXVlanRdData    <= "000000000000" & axiClkRXVlanRdData_i when (Bus2IP_RdCE(18) = '1') else (others => '0');
    axiClkRXVlanWrData_i  <= Bus2IP_Data(30 to 31);
    RxClClkRXVlanRdData   <= "000000000000" & rxClClkRxRdData_i;
  end generate RX_VLAN_STRP_TAG;

  RX_VLAN_STRP : if (C_RXVLAN_TRAN = 0 and C_RXVLAN_STRP = 1 and C_RXVLAN_TAG = 0) generate
  begin
    axiClkRXVlanRdData    <= "000000000000" & axiClkRXVlanRdData_i & '0' when (Bus2IP_RdCE(18) = '1') else (others => '0');
    axiClkRXVlanWrData_i  <= Bus2IP_Data(30 to 30);
    RxClClkRXVlanRdData   <= "000000000000" & rxClClkRxRdData_i & '0';
  end generate RX_VLAN_STRP;

  RX_VLAN_TAG : if (C_RXVLAN_TRAN = 0 and C_RXVLAN_STRP = 0 and C_RXVLAN_TAG = 1) generate
  begin
    axiClkRXVlanRdData    <= "000000000000" & '0' & axiClkRXVlanRdData_i when (Bus2IP_RdCE(18) = '1') else (others => '0');
    axiClkRXVlanWrData_i  <= Bus2IP_Data(31 to 31);
    RxClClkRXVlanRdData   <= "000000000000" & '0' & rxClClkRxRdData_i;
  end generate RX_VLAN_TAG;

  RX_VLAN_NONE : if (C_RXVLAN_TRAN = 0 and C_RXVLAN_STRP = 0 and C_RXVLAN_TAG = 0) generate
  begin
    axiClkRXVlanRdData    <= (others => '0');
    RxClClkRXVlanRdData   <= (others => '0');
  end generate RX_VLAN_NONE;

  IsRegData    <= isRegData_i;
  IeRegData    <= ieRegData_i;
  TtagRegData  <= ttagRegData_i;
  RtagRegData  <= rtagRegData_i;
  Tpid0RegData <= tpid0RegData_i;
  Tpid1RegData <= tpid1RegData_i;
  UawLRegData  <= uawLRegData_i;
  UawURegData  <= uawURegData_i;

  CR_I : reg_cr
    port map
    (
     Clk      => AxiClk,                -- in

     RST      => AxiReset,              -- in
     RdCE     => Bus2IP_RdCE(0),        -- in
     WrCE     => Bus2IP_WrCE(0),        -- in
     DataIn   => Bus2IP_Data(17 to 31), -- in
     DataOut  => crRdData,              -- out
     RegData  => CrRegData              -- out
    );

  TP_I : reg_tp
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(1),  -- in
     WrCE     => Bus2IP_WrCE(1),  -- in
     DataIn   => Bus2IP_Data(16 to 31), -- in
     DataOut  => tpRdData,          -- out
     RegData  => TpRegData,         -- out
     TPReq    => TPReq            -- out
    );

  IFGP_I : reg_ifgp
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(2),  -- in
     WrCE     => Bus2IP_WrCE(2),  -- in
     DataIn   => Bus2IP_Data(24 to 31), -- in
     DataOut  => ifgpRdData,          -- out
     RegData  => IfgpRegData          -- out
    );

  IS_I : reg_is
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(3),  -- in
     WrCE     => Bus2IP_WrCE(3),  -- in
     Intrpts  => IntrptsIn,         -- in
     DataIn   => Bus2IP_Data(23 to 31), -- out
     DataOut  => isRdData,          -- out
     RegData  => isRegData_i          -- out
    );

  IP_I : reg_ip
    port map
    (
     Clk      => AxiClk,              -- in
     RST      => AxiReset,      -- in
     RdCE     => Bus2IP_RdCE(4),    -- in
     IsIn     => isRegData_i,     -- in
     IeIn     => ieRegData_i,     -- in
     DataOut  => ipRdData,      -- out
     RegData  => IpRegData,     -- out
     Intrpt   => IntrptOut      -- out
    );

  IE_I : reg_ie
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(5),  -- in
     WrCE     => Bus2IP_WrCE(5),  -- in
     DataIn   => Bus2IP_Data(23 to 31), -- in
     DataOut  => ieRdData,          -- out
     RegData  => ieRegData_i          -- out
    );

  TTAG_I : reg_32b
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(6),  -- in
     WrCE     => Bus2IP_WrCE(6),  -- in
     DataIn   => Bus2IP_Data(0 to 31),  -- in
     DataOut  => ttagRdData,          -- out
     RegData  => ttagRegData_i          -- out
    );

  RTAG_I : reg_32b
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(7),  -- in
     WrCE     => Bus2IP_WrCE(7),  -- in
     DataIn   => Bus2IP_Data(0 to 31),  -- in
     DataOut  => rtagRdData,          -- out
     RegData  => rtagRegData_i          -- out
    );

  UAWL_I : reg_32b
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(8),  -- in
     WrCE     => Bus2IP_WrCE(8),  -- in
     DataIn   => Bus2IP_Data(0 to 31),  -- in
     DataOut  => uawLRdData,          -- out
     RegData  => uawLRegData_i         -- out
    );

  UAWU_I : reg_16bl
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(9),  -- in
     WrCE     => Bus2IP_WrCE(9),  -- in
     DataIn   => Bus2IP_Data(16 to 31), -- in
     DataOut  => uawURdData,          -- out
     RegData  => uawURegData_i          -- out
    );

  TPID0_I : reg_32b
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(10), -- in
     WrCE     => Bus2IP_WrCE(10), -- in
     DataIn   => Bus2IP_Data(0 to 31),  -- in
     DataOut  => tpid0RdData,         -- out
     RegData  => tpid0RegData_i        -- out
    );

  TPID1_I : reg_32b
    port map
    (
     Clk      => AxiClk,                  -- in
     RST      => AxiReset,          -- in
     RdCE     => Bus2IP_RdCE(11), -- in
     WrCE     => Bus2IP_WrCE(11), -- in
     DataIn   => Bus2IP_Data(0 to 31),  -- in
     DataOut  => tpid1RdData,         -- out
     RegData  => tpid1RegData_i        -- out
    );


  pcspma_status <= pcspma_status_cross when Bus2IP_RdCE(12) = '1' else (others => '0');


  EXTENDED_MULTICAST : if (C_MCAST_EXTEND = 1) generate
  begin

I_MULTICAST_MEM: xpm_memory_tdpram
  generic map (

    -- Common module generics
    MEMORY_SIZE             => 32768,            --positive integer
    MEMORY_PRIMITIVE        => "block",          --string; "auto", "distributed", "block" or "ultra" ;
    CLOCKING_MODE           => "independent_clock",  --string; "common_clock", "independent_clock" 
    MEMORY_INIT_FILE        => "none",          --string; "none" or "<filename>.mem" 
    MEMORY_INIT_PARAM       => "",              --string;
    USE_MEM_INIT            => 1,               --integer; 0,1
    WAKEUP_TIME             => "disable_sleep", --string; "disable_sleep" or "use_sleep_pin" 
    MESSAGE_CONTROL         => 0,               --integer;
    ECC_MODE                => "no_ecc",        --string; "no_ecc", "encode_only", "decode_only" or "both_encode_and_decode" 
    AUTO_SLEEP_TIME         => 0,               --Do not Change
    USE_EMBEDDED_CONSTRAINT => 0,               --integer: 0,1
    MEMORY_OPTIMIZATION     => "true",          --string; "true", "false" 

    -- Port A module generics
    WRITE_DATA_WIDTH_A      => 1,              --positive integer
    READ_DATA_WIDTH_A       => 1,              --positive integer
    BYTE_WRITE_WIDTH_A      => 1,              --integer; 8, 9, or WRITE_DATA_WIDTH_A value
    ADDR_WIDTH_A            => 15,               --positive integer
    READ_RESET_VALUE_A      => "0",             --string
    READ_LATENCY_A          => 1,               --non-negative integer
    WRITE_MODE_A            => "no_change",     --string; "write_first", "read_first", "no_change" 

    -- Port B module generics
    WRITE_DATA_WIDTH_B      => 1,              --positive integer
    READ_DATA_WIDTH_B       => 1,              --positive integer
    BYTE_WRITE_WIDTH_B      => 1,              --integer; 8, 9, or WRITE_DATA_WIDTH_B value
    ADDR_WIDTH_B            => 15,               --positive integer
    READ_RESET_VALUE_B      => "0",             --string
    READ_LATENCY_B          => 1,               --non-negative integer
    WRITE_MODE_B            => "no_change"      --string; "write_first", "read_first", "no_change" 
  )
  port map (

    -- Common module ports
    sleep                   => '0',

    -- Port A module ports
    clka                    => RxClClk,
    rsta                    => '0',
    ena                     => RxClClkMcastEn,
    regcea                  => '0',
    wea                     => "0",
    addra                   => RxClClkMcastAddr,
    dina                    => "0",
    injectsbiterra          => '0',
    injectdbiterra          => '0',
    douta                   => RxClClkMcastRdData,
    sbiterra                => open,
    dbiterra                => open,

    -- Port B module ports
    clkb                    => AxiClk,
    rstb                    => '0',
    enb                     => bus2IP_WrCE_20_en,
    regceb                  => '0',
    web                     => Bus2IP_WrCE(20 to 20),
    addrb                   => Bus2IP_Addr(15 to 29),
    dinb                    => Bus2IP_Data(31 to 31),
    injectsbiterrb          => '0',
    injectdbiterrb          => '0',
    doutb                   => AxiClkMcastRdData_i,
    sbiterrb                => open,
    dbiterrb                => open
  );

-- End of xpm_memory_tdpram_inst instance declaration

--    I_MULTICAST_MEM : entity lib_bmg_v1_0.blk_mem_gen_wrapper
--      generic map(
--        c_family                 => C_FAMILY,
--        c_xdevicefamily          => C_FAMILY,
--
--        -- Selection between BMG and XPM
--        bmg_xpm_sel              => 0,
--        -- Memory Specific Configurations
--        c_mem_type               => 2,
--           -- This wrapper only supports the True Dual Port RAM
--           -- 0: Single Port RAM
--           -- 1: Simple Dual Port RAM
--           -- 2: True Dual Port RAM
--           -- 3: Single Port Rom
--           -- 4: Dual Port RAM
--        c_algorithm              => 1,
--           -- 0: Selectable Primative
--           -- 1: Minimum Area
--        c_prim_type              => 0,
--           -- 0: ( 1-bit wide)
--           -- 1: ( 2-bit wide)
--           -- 2: ( 4-bit wide)
--           -- 3: ( 9-bit wide)
--           -- 4: (18-bit wide)
--           -- 5: (36-bit wide)
--           -- 6: (72-bit wide, single port only)
--        c_byte_size              => 8,   -- 8 or 9
--
--        -- Simulation Behavior Options
--        c_sim_collision_check    => "NONE",
--           -- "None"
--           -- "Generate_X"
--           -- "All"
--           -- "Warnings_only"
--        c_common_clk             => 0,   -- 0, 1
--        c_disable_warn_bhv_coll  => 0,   -- 0, 1
--        c_disable_warn_bhv_range => 0,   -- 0, 1
--
--        -- Initialization Configuration Options
--        c_load_init_file         => 0,
--        c_init_file_name         => "none",
--        c_use_default_data       => 0,   -- 0, 1
--        c_default_data           => "0", -- "..."
--
--        -- Port A Specific Configurations
--        c_has_mem_output_regs_a  => 0,   -- 0, 1
--        c_has_mux_output_regs_a  => 0,   -- 0, 1
--        c_write_width_a          => 1,  -- 1 to 1152
--        c_read_width_a           => 1,  -- 1 to 1152
--        c_write_depth_a          => 32768,  -- 2 to 9011200
--        c_read_depth_a           => 32768,  -- 2 to 9011200
--        c_addra_width            => 15,   -- 1 to 24
--        c_write_mode_a           => "NO_CHANGE",
--           -- "Write_First"
--           -- "Read_first"
--           -- "No_Change"
--        c_has_ena                => 1,   -- 0, 1
--        c_has_regcea             => 0,   -- 0, 1
--        c_has_ssra               => 0,   -- 0, 1
--        c_sinita_val             => "0", --"..."
--        c_use_byte_wea           => 0,   -- 0, 1
--        c_wea_width              => 1,   -- 1 to 128
--
--        -- Port B Specific Configurations
--        c_has_mem_output_regs_b  => 0,   -- 0, 1
--        c_has_mux_output_regs_b  => 0,   -- 0, 1
--        c_write_width_b          => 1,  -- 1 to 1152
--        c_read_width_b           => 1,  -- 1 to 1152
--        c_write_depth_b          => 32768,  -- 2 to 9011200
--        c_read_depth_b           => 32768,   -- 2 to 9011200
--        c_addrb_width            => 15,   -- 1 to 24
--        c_write_mode_b           => "NO_CHANGE",
--           -- "Write_First"
--           -- "Read_first"
--           -- "No_Change"
--        c_has_enb                => 0,   -- 0, 1
--        c_has_regceb             => 0,   -- 0, 1
--        c_has_ssrb               => 0,   -- 0, 1
--        c_sinitb_val             => "0", -- "..."
--        c_use_byte_web           => 0,   -- 0, 1
--        c_web_width              => 1,   -- 1 to 128
--
--        -- Other Miscellaneous Configurations
--        c_mux_pipeline_stages    => 0,   -- 0, 1, 2, 3
--           -- The number of pipeline stages within the MUX
--           --    for both Port A and Port B
--        c_use_ecc                => 0,
--           -- See DS512 for the limited core option selections for ECC support
--        c_use_ramb16bwer_rst_bhv => 0    --0, 1
--        )
--      port map
--        (
--        clka    => RxClClk,       --: in  std_logic;
--        ssra    => '0',            --: in  std_logic := '0';
--        dina    => "0",            --: in  std_logic_vector(c_write_width_a-1 downto 0) := (OTHERS => '0');
--        addra   => RxClClkMcastAddr,   --: in  std_logic_vector(c_addra_width-1   downto 0);
--        ena     => RxClClkMcastEn,     --: in  std_logic := '1';
--        regcea  => '0',            --: in  std_logic := '1';
--        wea     => "0",            --: in  std_logic_vector(c_wea_width-1     downto 0) := (OTHERS => '0');
--        douta   => RxClClkMcastRdData, --: out std_logic_vector(c_read_width_a-1  downto 0);
--
--        clkb    => AxiClk,    --: in  std_logic := '0';
--        ssrb    => '0',            --: in  std_logic := '0';
--        dinb    => Bus2IP_Data(31 to 31),--: in  std_logic_vector(c_write_width_b-1 downto 0) := (OTHERS => '0');
--        addrb   => Bus2IP_Addr(15 to 29),--: in  std_logic_vector(c_addrb_width-1   downto 0) := (OTHERS => '0');
--        enb     => bus2IP_WrCE_20_en,            --: in  std_logic := '1';
--        regceb  => '0',            --: in  std_logic := '1';
--        web     => Bus2IP_WrCE(20 to 20),--: in  std_logic_vector(c_web_width-1     downto 0) := (OTHERS => '0');
--        doutb   => AxiClkMcastRdData_i,--: out std_logic_vector(c_read_width_b-1  downto 0);
--
--        dbiterr => open,           --: out std_logic;
--           -- Double bit error that that cannot be auto corrected by ECC
--        sbiterr => open            --: out std_logic
--           -- Single Bit Error that has been auto corrected on the output bus
--        );
    AxiClkMcastRdData(0) <= AxiClkMcastRdData_i(0) and Bus2IP_RdCE(20);
  end generate EXTENDED_MULTICAST;

  NO_EXTENDED_MULTICAST : if (C_MCAST_EXTEND = 0) generate
  begin
    RxClClkMcastRdData <= (others => '0');
    AxiClkMcastRdData  <= (others => '0');
  end generate NO_EXTENDED_MULTICAST;

  TX_VLAN_BRAM : if (C_TXVLAN_TRAN = 1 or C_TXVLAN_TAG = 1 or C_TXVLAN_STRP = 1) generate
  begin

I_TX_VLAN_MEM: xpm_memory_tdpram
  generic map (

    -- Common module generics
    MEMORY_SIZE             => C_TXVLAN_WIDTH*4096,            --positive integer
    MEMORY_PRIMITIVE        => "block",          --string; "auto", "distributed", "block" or "ultra" ;
    CLOCKING_MODE           => "independent_clock",  --string; "common_clock", "independent_clock" 
    MEMORY_INIT_FILE        => "none",          --string; "none" or "<filename>.mem" 
    MEMORY_INIT_PARAM       => "",              --string;
    USE_MEM_INIT            => 1,               --integer; 0,1
    WAKEUP_TIME             => "disable_sleep", --string; "disable_sleep" or "use_sleep_pin" 
    MESSAGE_CONTROL         => 0,               --integer;
    ECC_MODE                => "no_ecc",        --string; "no_ecc", "encode_only", "decode_only" or "both_encode_and_decode" 
    AUTO_SLEEP_TIME         => 0,               --Do not Change
    USE_EMBEDDED_CONSTRAINT => 0,               --integer: 0,1
    MEMORY_OPTIMIZATION     => "true",          --string; "true", "false" 

    -- Port A module generics
    WRITE_DATA_WIDTH_A      => C_TXVLAN_WIDTH,              --positive integer
    READ_DATA_WIDTH_A       => C_TXVLAN_WIDTH,              --positive integer
    BYTE_WRITE_WIDTH_A      => C_TXVLAN_WIDTH,              --integer; 8, 9, or WRITE_DATA_WIDTH_A value
    ADDR_WIDTH_A            => 12,               --positive integer
    READ_RESET_VALUE_A      => "0",             --string
    READ_LATENCY_A          => 1,               --non-negative integer
    WRITE_MODE_A            => "no_change",     --string; "write_first", "read_first", "no_change" 

    -- Port B module generics
    WRITE_DATA_WIDTH_B      => C_TXVLAN_WIDTH,              --positive integer
    READ_DATA_WIDTH_B       => C_TXVLAN_WIDTH,              --positive integer
    BYTE_WRITE_WIDTH_B      => C_TXVLAN_WIDTH,              --integer; 8, 9, or WRITE_DATA_WIDTH_B value
    ADDR_WIDTH_B            => 12,               --positive integer
    READ_RESET_VALUE_B      => "0",             --string
    READ_LATENCY_B          => 1,               --non-negative integer
    WRITE_MODE_B            => "no_change"      --string; "write_first", "read_first", "no_change" 
  )
  port map (

    -- Common module ports
    sleep                   => '0',

    -- Port A module ports
    clka                    => AXI_STR_TXD_ACLK,
    rsta                    => '0',
    ena                     => AxiStrTxDClkTxVlanBramEnA,
    regcea                  => '0',
    wea                     => "0",
    addra                   => AxiStrTxDClkTxVlanAddr,
    dina                    => txvlan_dina,
    injectsbiterra          => '0',
    injectdbiterra          => '0',
    douta                   => AxiStrTxDClkTxRdData_i,
    sbiterra                => open,
    dbiterra                => open,

    -- Port B module ports
    clkb                    => AxiClk,
    rstb                    => '0',
    enb                     => bus2IP_WrCE_17_en,
    regceb                  => '0',
    web                     => Bus2IP_WrCE(17 to 17),
    addrb                   => Bus2IP_Addr(18 to 29),
    dinb                    => axiClkTxVlanWrData_i,
    injectsbiterrb          => '0',
    injectdbiterrb          => '0',
    doutb                   => axiClkTxVlanRdData_i,
    sbiterrb                => open,
    dbiterrb                => open
  );

-- End of xpm_memory_tdpram_inst instance declaration


--    I_TX_VLAN_MEM : entity lib_bmg_v1_0.blk_mem_gen_wrapper
--      generic map(
--        c_family                 => C_FAMILY,
--        c_xdevicefamily          => C_FAMILY,
--
--        -- Selection between BMG and XPM
--        bmg_xpm_sel              => 0,
--        -- Memory Specific Configurations
--        c_mem_type               => 2,
--           -- This wrapper only supports the True Dual Port RAM
--           -- 0: Single Port RAM
--           -- 1: Simple Dual Port RAM
--           -- 2: True Dual Port RAM
--           -- 3: Single Port Rom
--           -- 4: Dual Port RAM
--        c_algorithm              => 1,
--           -- 0: Selectable Primative
--           -- 1: Minimum Area
--        c_prim_type              => 3,
--           -- 0: ( 1-bit wide)
--           -- 1: ( 2-bit wide)
--           -- 2: ( 4-bit wide)
--           -- 3: ( 9-bit wide)
--           -- 4: (18-bit wide)
--           -- 5: (36-bit wide)
--           -- 6: (72-bit wide, single port only)
--        c_byte_size              => 8,   -- 8 or 9
--
--        -- Simulation Behavior Options
--        c_sim_collision_check    => "NONE",
--           -- "None"
--           -- "Generate_X"
--           -- "All"
--           -- "Warnings_only"
--        c_common_clk             => 0,   -- 0, 1
--        c_disable_warn_bhv_coll  => 0,   -- 0, 1
--        c_disable_warn_bhv_range => 0,   -- 0, 1
--
--        -- Initialization Configuration Options
--        c_load_init_file         => 0,
--        c_init_file_name         => "none",
--        c_use_default_data       => 0,   -- 0, 1
--        c_default_data           => "0", -- "..."
--
--        -- Port A Specific Configurations
--        c_has_mem_output_regs_a  => 0,   -- 0, 1
--        c_has_mux_output_regs_a  => 0,   -- 0, 1
--        c_write_width_a          => C_TXVLAN_WIDTH,  -- 1 to 1152
--        c_read_width_a           => C_TXVLAN_WIDTH,  -- 1 to 1152
--        c_write_depth_a          => 4096,  -- 2 to 9011200
--        c_read_depth_a           => 4096,  -- 2 to 9011200
--        c_addra_width            => 12,   -- 1 to 24
--        c_write_mode_a           => "NO_CHANGE",
--           -- "Write_First"
--           -- "Read_first"
--           -- "No_Change"
--        c_has_ena                => 0,   -- 0, 1
--        c_has_regcea             => 0,   -- 0, 1
--        c_has_ssra               => 0,   -- 0, 1
--        c_sinita_val             => "0", --"..."
--        c_use_byte_wea           => 0,   -- 0, 1
--        c_wea_width              => 1,   -- 1 to 128
--
--        -- Port B Specific Configurations
--        c_has_mem_output_regs_b  => 0,   -- 0, 1
--        c_has_mux_output_regs_b  => 0,   -- 0, 1
--        c_write_width_b          => C_TXVLAN_WIDTH,  -- 1 to 1152
--        c_read_width_b           => C_TXVLAN_WIDTH,  -- 1 to 1152
--        c_write_depth_b          => 4096,  -- 2 to 9011200
--        c_read_depth_b           => 4096,   -- 2 to 9011200
--        c_addrb_width            => 12,   -- 1 to 24
--        c_write_mode_b           => "NO_CHANGE",
--           -- "Write_First"
--           -- "Read_first"
--           -- "No_Change"
--        c_has_enb                => 0,   -- 0, 1
--        c_has_regceb             => 0,   -- 0, 1
--        c_has_ssrb               => 0,   -- 0, 1
--        c_sinitb_val             => "0", -- "..."
--        c_use_byte_web           => 0,   -- 0, 1
--        c_web_width              => 1,   -- 1 to 128
--
--        -- Other Miscellaneous Configurations
--        c_mux_pipeline_stages    => 0,   -- 0, 1, 2, 3
--           -- The number of pipeline stages within the MUX
--           --    for both Port A and Port B
--        c_use_ecc                => 0,
--           -- See DS512 for the limited core option selections for ECC support
--        c_use_ramb16bwer_rst_bhv => 0    --0, 1
--        )
--      port map
--        (
--        clka    => AXI_STR_TXD_ACLK,     --: in  std_logic;
--        ssra    => '0',            --: in  std_logic := '0';
--        dina    => txvlan_dina, --: in  std_logic_vector(c_write_width_a-1 downto 0) := (OTHERS => '0');
--        addra   => AxiStrTxDClkTxVlanAddr,  --: in  std_logic_vector(c_addra_width-1   downto 0);
--        ena     => AxiStrTxDClkTxVlanBramEnA,            --: in  std_logic := '1';
--        regcea  => '0',            --: in  std_logic := '1';
--        wea     => "0",            --: in  std_logic_vector(c_wea_width-1     downto 0) := (OTHERS => '0');
--        douta   => AxiStrTxDClkTxRdData_i,--: out std_logic_vector(c_read_width_a-1  downto 0);
--
--        clkb    => AxiClk,    --: in  std_logic := '0';
--        ssrb    => '0',            --: in  std_logic := '0';
--        dinb    => axiClkTxVlanWrData_i,--: in  std_logic_vector(c_write_width_b-1 downto 0) := (OTHERS => '0');
--        addrb   => Bus2IP_Addr(18 to 29),--: in  std_logic_vector(c_addrb_width-1   downto 0) := (OTHERS => '0');
--        enb     => bus2IP_WrCE_17_en,            --: in  std_logic := '1';
--        regceb  => '0',            --: in  std_logic := '1';
--        web     => Bus2IP_WrCE(17 to 17),--: in  std_logic_vector(c_web_width-1     downto 0) := (OTHERS => '0');
--        doutb   => axiClkTxVlanRdData_i,--: out std_logic_vector(c_read_width_b-1  downto 0);
--
--        dbiterr => open,           --: out std_logic;
--           -- Double bit error that that cannot be auto corrected by ECC
--        sbiterr => open            --: out std_logic
--           -- Single Bit Error that has been auto corrected on the output bus
--        );
  end generate TX_VLAN_BRAM;

  RX_VLAN_BRAM : if (C_RXVLAN_TRAN = 1 or C_RXVLAN_TAG = 1 or C_RXVLAN_STRP = 1) generate
  begin

I_RX_VLAN_MEM: xpm_memory_tdpram
  generic map (

    -- Common module generics
    MEMORY_SIZE             => C_RXVLAN_WIDTH*4096,            --positive integer
    MEMORY_PRIMITIVE        => "block",          --string; "auto", "distributed", "block" or "ultra" ;
    CLOCKING_MODE           => "independent_clock",  --string; "common_clock", "independent_clock" 
    MEMORY_INIT_FILE        => "none",          --string; "none" or "<filename>.mem" 
    MEMORY_INIT_PARAM       => "",              --string;
    USE_MEM_INIT            => 1,               --integer; 0,1
    WAKEUP_TIME             => "disable_sleep", --string; "disable_sleep" or "use_sleep_pin" 
    MESSAGE_CONTROL         => 0,               --integer;
    ECC_MODE                => "no_ecc",        --string; "no_ecc", "encode_only", "decode_only" or "both_encode_and_decode" 
    AUTO_SLEEP_TIME         => 0,               --Do not Change
    USE_EMBEDDED_CONSTRAINT => 0,               --integer: 0,1
    MEMORY_OPTIMIZATION     => "true",          --string; "true", "false" 

    -- Port A module generics
    WRITE_DATA_WIDTH_A      => C_RXVLAN_WIDTH,              --positive integer
    READ_DATA_WIDTH_A       => C_RXVLAN_WIDTH,              --positive integer
    BYTE_WRITE_WIDTH_A      => C_RXVLAN_WIDTH,              --integer; 8, 9, or WRITE_DATA_WIDTH_A value
    ADDR_WIDTH_A            => 12,               --positive integer
    READ_RESET_VALUE_A      => "0",             --string
    READ_LATENCY_A          => 1,               --non-negative integer
    WRITE_MODE_A            => "no_change",     --string; "write_first", "read_first", "no_change" 

    -- Port B module generics
    WRITE_DATA_WIDTH_B      => C_RXVLAN_WIDTH,              --positive integer
    READ_DATA_WIDTH_B       => C_RXVLAN_WIDTH,              --positive integer
    BYTE_WRITE_WIDTH_B      => C_RXVLAN_WIDTH,              --integer; 8, 9, or WRITE_DATA_WIDTH_B value
    ADDR_WIDTH_B            => 12,               --positive integer
    READ_RESET_VALUE_B      => "0",             --string
    READ_LATENCY_B          => 1,               --non-negative integer
    WRITE_MODE_B            => "no_change"      --string; "write_first", "read_first", "no_change" 
  )
  port map (

    -- Common module ports
    sleep                   => '0',

    -- Port A module ports
    clka                    => RxClClk,
    rsta                    => '0',
    ena                     => RxClClkRxVlanBramEnA,
    regcea                  => '0',
    wea                     => "0",
    addra                   => RxClClkRxVlanAddr,
    dina                    => rxvlan_dina,
    injectsbiterra          => '0',
    injectdbiterra          => '0',
    douta                   => rxClClkRxRdData_i,
    sbiterra                => open,
    dbiterra                => open,

    -- Port B module ports
    clkb                    => AxiClk,
    rstb                    => '0',
    enb                     => bus2IP_WrCE_18_en,
    regceb                  => '0',
    web                     => Bus2IP_WrCE(18 to 18),
    addrb                   => Bus2IP_Addr(18 to 29),
    dinb                    => axiClkRXVlanWrData_i,
    injectsbiterrb          => '0',
    injectdbiterrb          => '0',
    doutb                   => axiClkRXVlanRdData_i,
    sbiterrb                => open,
    dbiterrb                => open
  );

-- End of xpm_memory_tdpram_inst instance declaration


--    I_RX_VLAN_MEM : entity lib_bmg_v1_0.blk_mem_gen_wrapper
--      generic map(
--        c_family                 => C_FAMILY,
--        c_xdevicefamily          => C_FAMILY,
--
--        -- Selection between BMG and XPM
--        bmg_xpm_sel              => 0,
--        -- Memory Specific Configurations
--        c_mem_type               => 2,
--           -- This wrapper only supports the True Dual Port RAM
--           -- 0: Single Port RAM
--           -- 1: Simple Dual Port RAM
--           -- 2: True Dual Port RAM
--           -- 3: Single Port Rom
--           -- 4: Dual Port RAM
--        c_algorithm              => 1,
--           -- 0: Selectable Primative
--           -- 1: Minimum Area
--        c_prim_type              => 3,
--           -- 0: ( 1-bit wide)
--           -- 1: ( 2-bit wide)
--           -- 2: ( 4-bit wide)
--           -- 3: ( 9-bit wide)
--           -- 4: (18-bit wide)
--           -- 5: (36-bit wide)
--           -- 6: (72-bit wide, single port only)
--        c_byte_size              => 8,   -- 8 or 9
--
--        -- Simulation Behavior Options
--        c_sim_collision_check    => "NONE",
--           -- "None"
--           -- "Generate_X"
--           -- "All"
--           -- "Warnings_only"
--        c_common_clk             => 0,   -- 0, 1
--        c_disable_warn_bhv_coll  => 0,   -- 0, 1
--        c_disable_warn_bhv_range => 0,   -- 0, 1
--
--        -- Initialization Configuration Options
--        c_load_init_file         => 0,
--        c_init_file_name         => "none",
--        c_use_default_data       => 0,   -- 0, 1
--        c_default_data           => "0", -- "..."
--
--        -- Port A Specific Configurations
--        c_has_mem_output_regs_a  => 0,   -- 0, 1
--        c_has_mux_output_regs_a  => 0,   -- 0, 1
--        c_write_width_a          => C_RXVLAN_WIDTH,  -- 1 to 1152
--        c_read_width_a           => C_RXVLAN_WIDTH,  -- 1 to 1152
--        c_write_depth_a          => 4096,  -- 2 to 9011200
--        c_read_depth_a           => 4096,  -- 2 to 9011200
--        c_addra_width            => 12,   -- 1 to 24
--        c_write_mode_a           => "NO_CHANGE",
--           -- "Write_First"
--           -- "Read_first"
--           -- "No_Change"
--        c_has_ena                => 0,   -- 0, 1
--        c_has_regcea             => 0,   -- 0, 1
--        c_has_ssra               => 0,   -- 0, 1
--        c_sinita_val             => "0", --"..."
--        c_use_byte_wea           => 0,   -- 0, 1
--        c_wea_width              => 1,   -- 1 to 128
--
--        -- Port B Specific Configurations
--        c_has_mem_output_regs_b  => 0,   -- 0, 1
--        c_has_mux_output_regs_b  => 0,   -- 0, 1
--        c_write_width_b          => C_RXVLAN_WIDTH,  -- 1 to 1152
--        c_read_width_b           => C_RXVLAN_WIDTH,  -- 1 to 1152
--        c_write_depth_b          => 4096,  -- 2 to 9011200
--        c_read_depth_b           => 4096,   -- 2 to 9011200
--        c_addrb_width            => 12,   -- 1 to 24
--        c_write_mode_b           => "NO_CHANGE",
--           -- "Write_First"
--           -- "Read_first"
--           -- "No_Change"
--        c_has_enb                => 0,   -- 0, 1
--        c_has_regceb             => 0,   -- 0, 1
--        c_has_ssrb               => 0,   -- 0, 1
--        c_sinitb_val             => "0", -- "..."
--        c_use_byte_web           => 0,   -- 0, 1
--        c_web_width              => 1,   -- 1 to 128
--
--        -- Other Miscellaneous Configurations
--        c_mux_pipeline_stages    => 0,   -- 0, 1, 2, 3
--           -- The number of pipeline stages within the MUX
--           --    for both Port A and Port B
--        c_use_ecc                => 0,
--           -- See DS512 for the limited core option selections for ECC support
--        c_use_ramb16bwer_rst_bhv => 0    --0, 1
--        )
--      port map
--        (
--        clka    => RxClClk,     --: in  std_logic;
--        ssra    => '0',            --: in  std_logic := '0';
--        dina    => rxvlan_dina, --: in  std_logic_vector(c_write_width_a-1 downto 0) := (OTHERS => '0');
--        addra   => RxClClkRxVlanAddr,  --: in  std_logic_vector(c_addra_width-1   downto 0);
--        ena     => RxClClkRxVlanBramEnA,            --: in  std_logic := '1';
--        regcea  => '0',            --: in  std_logic := '1';
--        wea     => "0",            --: in  std_logic_vector(c_wea_width-1     downto 0) := (OTHERS => '0');
--        douta   => rxClClkRxRdData_i,--: out std_logic_vector(c_read_width_a-1  downto 0);
--
--        clkb    => AxiClk,    --: in  std_logic := '0';
--        ssrb    => '0',            --: in  std_logic := '0';
--        dinb    => axiClkRXVlanWrData_i,--: in  std_logic_vector(c_write_width_b-1 downto 0) := (OTHERS => '0');
--        addrb   => Bus2IP_Addr(18 to 29),--: in  std_logic_vector(c_addrb_width-1   downto 0) := (OTHERS => '0');
--        enb     => bus2IP_WrCE_18_en,            --: in  std_logic := '1';
--        regceb  => '0',            --: in  std_logic := '1';
--        web     => Bus2IP_WrCE(18 to 18),--: in  std_logic_vector(c_web_width-1     downto 0) := (OTHERS => '0');
--        doutb   => axiClkRXVlanRdData_i,--: out std_logic_vector(c_read_width_b-1  downto 0);
--
--        dbiterr => open,           --: out std_logic;
--           -- Double bit error that that cannot be auto corrected by ECC
--        sbiterr => open            --: out std_logic
--           -- Single Bit Error that has been auto corrected on the output bus
--        );
  end generate RX_VLAN_BRAM;

  RD_ACK_BLOCKER_PROCESS : process (AxiClk,AxiReset)
  begin
    if (AxiClk'event and AxiClk = '1') then
      if (AxiReset = '1') then
        rdAckBlocker <= '0';
      else
        rdAckBlocker <= (softRead_d1) or  -- set when = '1'
                        (rdAckBlocker and -- hold  when = '1'
                        (softRead_d1));   -- clear when = '0'
      end if;
    end if;
  end process;

  WR_ACK_BLOCKER_PROCESS : process (AxiClk,AxiReset)
  begin
    if (AxiClk'event and AxiClk = '1') then
      if (AxiReset = '1') then
        wrAckBlocker <= '0';
      else
        wrAckBlocker <= (softWrite_d1) or -- set when = '1'
                        (wrAckBlocker and -- hold  when = '1'
                        (softWrite_d1));  -- clear when = '0'
      end if;
    end if;
  end process;

  --------------------------------------------------------------------------
  -- ACK_PROCESS
  --------------------------------------------------------------------------
  ACK_PROCESS : process (AxiReset, AxiClk)
  begin
    if (AxiClk'event and AxiClk = '1') then
      if (AxiReset = '1') then
        softRead_d1  <= '0';
        softWrite_d1 <= '0';
        iP2Bus_WrAck_i  <= '0';
        iP2Bus_RdAck_i  <= '0';
      else
        softRead_d1  <= softRead;
        softWrite_d1 <= softWrite;
        iP2Bus_WrAck_i  <= ( softWrite_d1) and not(wrAckBlocker);
        iP2Bus_RdAck_i  <= ( softRead_d1) and not(rdAckBlocker);
      end if;
    end if;
  end process;

  softRead    <= Bus2IP_RdCE(0) or
                 Bus2IP_RdCE(1) or
                 Bus2IP_RdCE(2) or
                 Bus2IP_RdCE(3) or
                 Bus2IP_RdCE(4) or
                 Bus2IP_RdCE(5) or
                 Bus2IP_RdCE(6) or
                 Bus2IP_RdCE(7) or
                 Bus2IP_RdCE(8) or
                 Bus2IP_RdCE(9) or
                 Bus2IP_RdCE(10) or
                 Bus2IP_RdCE(11) or
                 Bus2IP_RdCE(12) or
                 Bus2IP_RdCE(17) or
                 Bus2IP_RdCE(18) or
                 Bus2IP_RdCE(20);
  softWrite   <= Bus2IP_WrCE(0) or
                 Bus2IP_WrCE(1) or
                 Bus2IP_WrCE(2) or
                 Bus2IP_WrCE(3) or
                 Bus2IP_WrCE(4) or
                 Bus2IP_WrCE(5) or
                 Bus2IP_WrCE(6) or
                 Bus2IP_WrCE(7) or
                 Bus2IP_WrCE(8) or
                 Bus2IP_WrCE(9) or
                 Bus2IP_WrCE(10) or
                 Bus2IP_WrCE(11) or
                 Bus2IP_WrCE(17) or
                 Bus2IP_WrCE(18) or
                 Bus2IP_WrCE(20);

  rdData  <= (
              ("00000000000000000" & crRdData) or
              ("0000000000000000" & tpRdData) or
              ("000000000000000000000000" & ifgpRdData)or
              ("00000000000000000000000" & isRdData) or
              ("00000000000000000000000" & ieRdData) or
              ("00000000000000000000000" & ipRdData) or
              ttagRdData or
              rtagRdData or
              tpid0RdData or
              tpid1RdData or
              ("0000000000000000" & pcspma_status) or
              uawLRdData or
              ("0000000000000000" & uawURdData) or
              ("0000000000000000000000000000000" & AxiClkMcastRdData) or
              ("000000000000000000" & axiClkTxVlanRdData) or
              ("000000000000000000" & axiClkRXVlanRdData)
             );

  --------------------------------------------------------------------------
  -- ACK_RD_DATA_PROCESS
  --------------------------------------------------------------------------
  ACK_RD_DATA_PROCESS : process (AxiReset, AxiClk)
  begin
    if (AxiClk'event and AxiClk = '1') then
      if (AxiReset = '1') then
        IP2Bus_WrAck <= '0';
        IP2Bus_RdAck <= '0';
        IP2Bus_Data  <= (others => '0');
      else
        IP2Bus_WrAck <= iP2Bus_WrAck_i;
        IP2Bus_RdAck <= iP2Bus_RdAck_i;
        IP2Bus_Data  <= rdData;
      end if;
    end if;
  end process;

end imp;


------------------------------------------------------------------------
-- Title      : Package for the tri_mode_ethernet_fifo logic
-- Project    : Tri-Mode Ethernet FIFO
------------------------------------------------------------------------
-- File       : axi_ethernet_buffer_v2_0_25_pack.vhd
-- Author     : Xilinx Inc.
------------------------------------------------------------------------
-- (c) Copyright 2012 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
------------------------------------------------------------------------
-- Description:  This package contains all component declarations for
--               the entiries which make up the Tx I/F logic
------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

library axi_lite_ipif_v3_0_5;
use axi_lite_ipif_v3_0_5.all;

package axi_ethernet_buffer_v2_0_25_pack is

  ----------------------------------------------------------------------------
  --  Component Declarations
  ----------------------------------------------------------------------------
  component reset_combiner
  generic (
    C_PHY_RST_COUNT       : integer   := 1321; 
    C_FAMILY               : string                        := "virtex7";
    C_SIMULATION         : integer range 0 to 1 := 0
  );
  port (
    S_AXI_ACLK           : in  std_logic;   --  AXI4-Lite Clock
    S_AXI_ARESETN        : in  std_logic;   --  AXI4-Lite Reset
    GTX_CLK_125MHZ       : in  std_logic;   --  GTX CLK
    RX_CLIENT_CLK        : in  std_logic;   --  Receive Client Clock
    RX_CLIENT_CLK_EN     : in  std_logic;   --  Receive Client Clock Enable
    TX_CLIENT_CLK        : in  std_logic;   --  Transmit Client Clock
    TX_CLIENT_CLK_EN     : in  std_logic;   --  Transmit Client Clock Enable
    AXI_STR_TXD_ACLK     : in  std_logic;   --  AXI-Stream Transmit Clock
    AXI_STR_TXD_ARESETN  : in  std_logic;   --  AXI-Stream Transmit Reset
    AXI_STR_TXC_ACLK     : in  std_logic;   --  AXI-Stream Transmit Clock
    AXI_STR_TXC_ARESETN  : in  std_logic;   --  AXI-Stream Transmit Reset
    AXI_STR_RXD_ACLK     : in  std_logic;   --  AXI-Stream Receive Clock
    AXI_STR_RXD_ARESETN  : in  std_logic;   --  AXI-Stream Receive Reset
    AXI_STR_RXS_ACLK     : in  std_logic;   --  AXI-Stream Receive Clock
    AXI_STR_RXS_ARESETN  : in  std_logic;   --  AXI-Stream Receive Reset
    PHY_RESET_N          : out std_logic;   --  PHY Reset
    PHY_RESET_CMPLTE     : out std_logic;   --  PHY Reset Complete
    RESET2AXI            : out std_logic;   --  Reset going to AXI
    RESET2RX_CLIENT      : out std_logic;   --  Reset going to Receive Client Interface
    RESET2TX_CLIENT      : out std_logic;   --  Reset going to Transmit Client Interface
    RESET2AXI_STR_TXD    : out std_logic;   --  Reset going to AXI-Stream Transmit Data Interface
    RESET2AXI_STR_TXC    : out std_logic;   --  Reset going to AXI-Stream Transmit Control Interface
    RESET2AXI_STR_RXD    : out std_logic;   --  Reset going to AXI-Stream Receive Data Interface
    RESET2AXI_STR_RXS    : out std_logic;   --  Reset going to AXI-Stream Receive Status Interface
    RESET2GTX_CLK        : out std_logic    --  Reset going to GTX Clock signals
  );
  end component;
  component addr_response_shim
  generic (

      C_BUS2CORE_CLK_RATIO      : integer range 1 to 2    := 1;
      C_S_AXI_ADDR_WIDTH        : integer range 32 to 32  := 32;
      C_S_AXI_DATA_WIDTH        : integer range 32 to 32  := 32;
      C_SIPIF_DWIDTH            : integer range 32 to 32  := 32;
      C_NUM_CS                  : integer                 := 10;
      C_NUM_CE                  : integer                 := 41;
      C_FAMILY                  : string                  := "virtex6"
      );
  port (
      --Clock and Reset
      BUS2IP_CLK                : in  std_logic;                                        --  AXI4-Lite clk
      BUS2IP_RESET              : in  std_logic;                                        --  AXI4-Lite reset

      -- PLB Slave Interface with Shim
      BUS2IP_ADDR             : in  std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );   --  Address bus from AXI4-Lite to Shim
      BUS2IP_DATA             : in  std_logic_vector(0 to C_SIPIF_DWIDTH - 1 );       --  Data bus from AXI4-Lite to Shim
      BUS2IP_RNW              : in  std_logic;                                        --  RNW signal from AXI4-Lite to Shim
      BUS2IP_CS               : in  std_logic_vector(0 to 0);                         --  CS signal from AXI4-Lite to Shim
      BUS2IP_RdCE             : in  std_logic_vector(0 to 0);                         --  RdCE signal from AXI4-Lite to Shim
      BUS2IP_WrCE             : in  std_logic_vector(0 to 0);                         --  WrCE signal from AXI4-Lite to Shim

      IP2BUS_DATA             : out std_logic_vector (0 to C_SIPIF_DWIDTH - 1 );      --  Data bus from Shim to AXI4-Lite
      IP2BUS_WrAck            : out std_logic;                                        --  WrCE signal from Shim to AXI4-Lite
      IP2BUS_RdAck            : out std_logic;                                        --  RdCE signal from Shim to AXI4-Lite

      -- TEMAC Interface with Shim
      Shim2IP_Addr              : out std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );   --  Address bus from Shim to AXI Ethernet
      Shim2IP_Data              : out std_logic_vector(0 to C_SIPIF_DWIDTH - 1 );       --  Data bus from Shim to AXI Ethernet
      Shim2IP_RNW               : out std_logic;                                        --  RNW signal from Shim to AXI Ethernet
      Shim2IP_CS                : out std_logic_vector(0 to C_NUM_CS);                  --  CS signal from Shim to AXI Ethernet
      Shim2IP_RdCE              : out std_logic_vector(0 to C_NUM_CE);                  --  RdCE signal from Shim to AXI Ethernet
      Shim2IP_WrCE              : out std_logic_vector(0 to C_NUM_CE);                  --  WrCE signal from Shim to AXI Ethernet

      IP2Shim_Data              : in  std_logic_vector (0 to C_SIPIF_DWIDTH - 1 );      --  Data bus from AXI Ethernet to Shim
      IP2Shim_WrAck             : in  std_logic;                                        --  WrCE signal from AXI Ethernet to Shim
      IP2Shim_RdAck             : in  std_logic                                         --  RdCE signal from AXI Ethernet to Shim
   );

  end component;
  component axi_ethernet_buffer_v2_0_25 
  generic (
    --  System Generics
    C_FAMILY               : string                        := "virtex7";
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32        := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32        := 32;
    C_TEMAC_ADDR_WIDTH     : integer range 0 to 32        := 12;
    C_HALFDUP              : integer range 0 to 1          := 0;
    C_TXMEM                : integer                       := 4096;
    C_ENABLE_1588       : integer    := 0;
    C_RXMEM                : integer                       := 4096;
    C_TXCSUM               : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_RXCSUM               : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_TXVLAN_TRAN          : integer range 0 to 1          := 0;
    C_RXVLAN_TRAN          : integer range 0 to 1          := 0;
    C_TXVLAN_TAG           : integer range 0 to 1          := 0;
    C_RXVLAN_TAG           : integer range 0 to 1          := 0;
    C_TXVLAN_STRP          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP          : integer range 0 to 1          := 0;
    C_MCAST_EXTEND         : integer range 0 to 1          := 0;
    C_SIMULATION           : integer                       := 0;

    C_AVB                 : integer range 0 to 1          := 0;
    C_STATS               : integer range 0 to 1          := 0;
    C_ENABLE_LVDS         : integer range 0 to 1          := 0;
    C_PHY_TYPE            : integer range 0 to 5          := 1;
    C_PHYADDR             : integer range 0 to 31    := 1; 
    C_PHY_RST_COUNT       : integer   := 1321; 
    C_TYPE                : integer range 0 to 2          := 0
  );
  port (
    -- System signals ---------------------------------------------------------
    S_AXI_ACLK              : in  std_logic;                                        
    S_AXI_ARESETN           : in  std_logic;                                        
    INTERRUPT               : out std_logic;                                        --  AXI Ethernet Interrupt
    -- AXI Lite signals
    S_AXI_AWADDR            : in  std_logic_vector (17 downto 0);
    S_AXI_AWVALID           : in  std_logic;                                        
    S_AXI_AWREADY           : out std_logic;                                        
    S_AXI_WDATA             : in  std_logic_vector  (31 downto 0);
    S_AXI_WSTRB             : in  std_logic_vector (3 downto 0);
    S_AXI_WVALID            : in  std_logic;                                        
    S_AXI_WREADY            : out std_logic;                                        
    S_AXI_BRESP             : out std_logic_vector(1 downto 0);                     
    S_AXI_BVALID            : out std_logic;                                        
    S_AXI_BREADY            : in  std_logic;                                        
    S_AXI_ARADDR            : in  std_logic_vector (17 downto 0);
    S_AXI_ARVALID           : in  std_logic;                                        
    S_AXI_ARREADY           : out std_logic;                                        
    S_AXI_RDATA             : out std_logic_vector (31 downto 0);
    S_AXI_RRESP             : out std_logic_vector(1 downto 0);                     
    S_AXI_RVALID            : out std_logic;                                        
    S_AXI_RREADY            : in  std_logic;                                        


    -- Interrupt sources
    EMAC_CLIENT_AUTONEG_INT : in  std_logic;                                        --  Auto negotiation signal from EMAC
    EMAC_RESET_DONE_INT     : in  std_logic;                                        --  Reset Done signal from EMAC
    EMAC_RX_DCM_LOCKED_INT  : in  std_logic;                                        --  DCM Locked signal from EMAC
    PCSPMA_STATUS_VECTOR    : in  std_logic_vector(15 downto 0);                    --  Link Status vector from PCS/PMA core
--    TEMAC_IPIC2GHI_INTR     : in  std_logic;                                        --  Interrupt


    -- AXI Stream signals
    AXI_STR_TXD_ACLK      : in  std_logic;                                          --  AXI-Stream Transmit Data Clk
    AXI_STR_TXD_ARESETN   : in  std_logic;                                          --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID    : in  std_logic;                                          --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY    : out std_logic;                                          --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST     : in  std_logic;                                          --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TKEEP     : in  std_logic_vector(3 downto 0);                       --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA     : in  std_logic_vector(31 downto 0);                      --  AXI-Stream Transmit Data Data

    AXI_STR_TXC_ACLK      : in  std_logic;                                          --  AXI-Stream Transmit Control Clk
    AXI_STR_TXC_ARESETN   : in  std_logic;                                          --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID    : in  std_logic;                                          --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY    : out std_logic;                                          --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST     : in  std_logic;                                          --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TKEEP     : in  std_logic_vector(3 downto 0);                       --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA     : in  std_logic_vector(31 downto 0);                      --  AXI-Stream Transmit Control Data

    AXI_STR_RXD_ACLK        : in  std_logic;                                        --  AXI-Stream Receive Data Clk
    AXI_STR_RXD_ARESETN     : in  std_logic;                                        --  AXI-Stream Receive Data Reset
    AXI_STR_RXD_VALID       : out std_logic;                                        --  AXI-Stream Receive Data Valid
    AXI_STR_RXD_READY       : in  std_logic;                                        --  AXI-Stream Receive Data Ready
    AXI_STR_RXD_LAST        : out std_logic;                                        --  AXI-Stream Receive Data Last
    AXI_STR_RXD_KEEP        : out std_logic_vector(3 downto 0);                     --  AXI-Stream Receive Data Keep
    AXI_STR_RXD_DATA        : out std_logic_vector(31 downto 0);                    --  AXI-Stream Receive Data Data

    AXI_STR_RXS_ACLK        : in  std_logic;                                        --  AXI-Stream Receive Status Clk
    AXI_STR_RXS_ARESETN     : in  std_logic;                                        --  AXI-Stream Receive Status Reset
    AXI_STR_RXS_VALID       : out std_logic;                                        --  AXI-Stream Receive Status Valid
    AXI_STR_RXS_READY       : in  std_logic;                                        --  AXI-Stream Receive Status Ready
    AXI_STR_RXS_LAST        : out std_logic;                                        --  AXI-Stream Receive Status Last
    AXI_STR_RXS_KEEP        : out std_logic_vector(3 downto 0);                     --  AXI-Stream Receive Status Keep
    AXI_STR_RXS_DATA        : out std_logic_vector(31 downto 0);                    --  AXI-Stream Receive Status Data

    -- TEMAC Interface
    ------------------------
    pause_req               : out std_logic;                                        -- pause req from register to TEMAC
    pause_val               : out std_logic_vector(16 to 31);                       -- pause value from register to TEMAC

  ------------------------------
    -- Signals added for axi lite split logic
    S_AXI_2TEMAC_AWADDR : out STD_LOGIC_VECTOR ( C_TEMAC_ADDR_WIDTH - 1 downto 0 );
    S_AXI_2TEMAC_AWVALID : out STD_LOGIC;
    S_AXI_2TEMAC_AWREADY : in STD_LOGIC;
    S_AXI_2TEMAC_WDATA : out STD_LOGIC_VECTOR ( 31 downto 0 );
    S_AXI_2TEMAC_WVALID : out STD_LOGIC;
    S_AXI_2TEMAC_WREADY : in STD_LOGIC;
    S_AXI_2TEMAC_BRESP : in STD_LOGIC_VECTOR ( 1 downto 0 );
    S_AXI_2TEMAC_BVALID : in STD_LOGIC;
    S_AXI_2TEMAC_BREADY : out STD_LOGIC;
    S_AXI_2TEMAC_ARADDR : out STD_LOGIC_VECTOR ( C_TEMAC_ADDR_WIDTH - 1 downto 0 );
    S_AXI_2TEMAC_ARVALID : out STD_LOGIC;
    S_AXI_2TEMAC_ARREADY : in STD_LOGIC;
    S_AXI_2TEMAC_RDATA : in STD_LOGIC_VECTOR ( 31 downto 0 );
    S_AXI_2TEMAC_RRESP : in STD_LOGIC_VECTOR ( 1 downto 0 );
    S_AXI_2TEMAC_RVALID : in STD_LOGIC;
    S_AXI_2TEMAC_RREADY : out STD_LOGIC;
    -- end of Signals added for axi lite split logic
  ------------------------------

    -- added 05/5/2011
    RX_CLK_ENABLE_IN        : in std_logic;                                         -- TEMAC clock domain enable

    rx_statistics_vector    : in  std_logic_vector(27 downto 0);                    -- RX statistics from TEMAC
    rx_statistics_valid     : in  std_logic;                                        -- Rx stats valid from TEMAC

    rx_mac_aclk             : in  std_logic;                                        -- Rx axistream clock from TEMAC
    rx_reset                : in  std_logic;                                        -- Rx axistream reset from TEMAC
    rx_axis_mac_tdata       : in  std_logic_vector(7 downto 0);                     -- Rx axistream data from TEMAC
    rx_axis_mac_tvalid      : in  std_logic;                                        -- Rx axistream valid from TEMAC
    rx_axis_mac_tlast       : in  std_logic;                                        -- Rx axistream last from TEMAC
    rx_axis_mac_tuser       : in  std_logic;                                        -- Rx axistream good/bad indicator from TEMAC

    tx_ifg_delay            : out std_logic_vector(24 to 31);                       -- interframe gap delay from register to TEMAC

    tx_mac_aclk             : in  std_logic;                                        -- Tx axistream clock from TEMAC
    tx_reset                : in  std_logic;                                        -- Tx axistream reset from TEMAC
    tx_axis_mac_tdata       : out std_logic_vector(7 downto 0);                     -- Tx axistream data to TEMAC
    tx_axis_mac_tvalid      : out std_logic;                                        -- Tx axistream valid to TEMAC
    tx_axis_mac_tlast       : out std_logic;                                        -- Tx axistream last to TEMAC
    tx_axis_mac_tuser       : out std_logic_vector(0 downto 0);                                        -- Tx axistream underrun indicator to TEMAC
    tx_axis_mac_tready      : in  std_logic;                                        -- Tx axistream ready from TEMAC
--    tx_collision            : in  std_logic;                                        -- Tx collision not used from TEMAC
--    tx_retransmit           : in  std_logic;                                        -- Tx retransmit not used from TEMAC

    speed_is_10_100         : in  std_logic;                                        -- speed is 10/100 not 1000 indicator

    RESET2PCSPMA                     : out std_logic;                                --  Reset to TEMAC
    RESET2TEMACn                    : out std_logic;                                --  Reset to TEMAC (active low version)

    -- Ethernet System signals -----------------------------------------------
    PHY_RST_N                       : out std_logic;                                --  Reset to PHY

    mdio_i_top          : in   std_logic; -- input from top
    mdio_o_top    : out  std_logic;
    mdio_t_top    : out  std_logic;
    mdc_top       : out  std_logic;
    mdio_t_pcspma       : in   std_logic; -- input from pcspma
    mdio_o_pcspma       : in   std_logic; -- input from pcspma
    mdio_i_temac  : out  std_logic; -- output to temac
    mdio_o_temac  : in   std_logic;
    mdio_t_temac  : in   std_logic;
    mdc_temac     : in   std_logic;

    -- GTX_CLK 125 MHz clock
    GTX_CLK                         : in  std_logic                                 --  GTX CLK


  );

  end component;
-----  component axi_ethernet_buffer_v2_0_25
-----  generic (
-----    --  System Generics
-----    C_FAMILY               : string                        := "virtex7";
-----    C_HAS_SGMII            : integer range 0 to 1          := 0;
-----    C_S_AXI_ACLK_FREQ_HZ   : INTEGER                       := 100000000;
-----    --  Frequency of the AXI clock in Hertz auto computed by the tools
-----    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32        := 32;
-----    C_S_AXI_DATA_WIDTH     : integer range 32 to 32        := 32;
-----    C_S_AXI_ID_WIDTH       : INTEGER range 1 to 4          := 4;
-----    C_HALFDUP              : integer range 0 to 1          := 0;
-----    C_TXMEM                : integer                       := 4096;
-----    C_RXMEM                : integer                       := 4096;
-----    C_TXCSUM               : integer range 0 to 2          := 0;
-----      -- 0 - No checksum offloading
-----      -- 1 - Partial (legacy) checksum offloading
-----      -- 2 - Full checksum offloading
-----    C_RXCSUM               : integer range 0 to 2          := 0;
-----      -- 0 - No checksum offloading
-----      -- 1 - Partial (legacy) checksum offloading
-----      -- 2 - Full checksum offloading
-----    C_TXVLAN_TRAN          : integer range 0 to 1          := 0;
-----    C_RXVLAN_TRAN          : integer range 0 to 1          := 0;
-----    C_TXVLAN_TAG           : integer range 0 to 1          := 0;
-----    C_RXVLAN_TAG           : integer range 0 to 1          := 0;
-----    C_TXVLAN_STRP          : integer range 0 to 1          := 0;
-----    C_RXVLAN_STRP          : integer range 0 to 1          := 0;
-----    C_MCAST_EXTEND         : integer range 0 to 1          := 0;
-----    C_SIMULATION           : integer                       := 0
-----  );
-----  port (
-----    -- IPIF control signals
-----    INTERRUPT               : out std_logic;                                        --  AXI Ethernet Interrupt
-----    BUS2IP_CLK              : in  std_logic;                                        --  AXI4-Lite Clk to top level
-----    BUS2IP_RESET            : in  std_logic;                                        --  AXI4-Lite Reset to top level
-----    BUS2IP_CS               : in  std_logic_vector(0 to 0);
-----    BUS2IP_RDCE             : in  std_logic_vector(0 to 0);
-----    BUS2IP_WRCE             : in  std_logic_vector(0 to 0);
-----    BUS2IP_ADDR             : in  std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );
-----    BUS2IP_DATA             : in  std_logic_vector(0 to C_S_AXI_DATA_WIDTH - 1 );
-----    BUS2IP_R_NW             : in  std_logic;
-----    IP2BUS_DATA             : out std_logic_vector (0 to C_S_AXI_DATA_WIDTH - 1 );
-----    IP2BUS_WR_ACK           : out std_logic;
-----    IP2BUS_RD_ACK           : out std_logic;
-----
-----    -- Interrupt sources
-----    EMAC_CLIENT_AUTONEG_INT : in  std_logic;                                        --  Auto negotiation signal from EMAC
-----    EMAC_RESET_DONE_INT     : in  std_logic;                                        --  Reset Done signal from EMAC
-----    EMAC_RX_DCM_LOCKED_INT  : in  std_logic;                                        --  DCM Locked signal from EMAC
-----    PCSPMA_STATUS_VECTOR    : in  std_logic_vector(15 downto 0);                    --  Link Status vector from PCS/PMA core
-----
-----
-----    -- AXI Stream signals
-----    AXI_STR_TXD_ACLK      : in  std_logic;                                          --  AXI-Stream Transmit Data Clk
-----    AXI_STR_TXD_ARESETN   : in  std_logic;                                          --  AXI-Stream Transmit Data Reset
-----    AXI_STR_TXD_TVALID    : in  std_logic;                                          --  AXI-Stream Transmit Data Valid
-----    AXI_STR_TXD_TREADY    : out std_logic;                                          --  AXI-Stream Transmit Data Ready
-----    AXI_STR_TXD_TLAST     : in  std_logic;                                          --  AXI-Stream Transmit Data Last
-----    AXI_STR_TXD_TKEEP     : in  std_logic_vector(3 downto 0);                       --  AXI-Stream Transmit Data Keep
-----    AXI_STR_TXD_TDATA     : in  std_logic_vector(31 downto 0);                      --  AXI-Stream Transmit Data Data
-----
-----    AXI_STR_TXC_ACLK      : in  std_logic;                                          --  AXI-Stream Transmit Control Clk
-----    AXI_STR_TXC_ARESETN   : in  std_logic;                                          --  AXI-Stream Transmit Control Reset
-----    AXI_STR_TXC_TVALID    : in  std_logic;                                          --  AXI-Stream Transmit Control Valid
-----    AXI_STR_TXC_TREADY    : out std_logic;                                          --  AXI-Stream Transmit Control Ready
-----    AXI_STR_TXC_TLAST     : in  std_logic;                                          --  AXI-Stream Transmit Control Last
-----    AXI_STR_TXC_TKEEP     : in  std_logic_vector(3 downto 0);                       --  AXI-Stream Transmit Control Keep
-----    AXI_STR_TXC_TDATA     : in  std_logic_vector(31 downto 0);                      --  AXI-Stream Transmit Control Data
-----
-----    AXI_STR_RXD_ACLK        : in  std_logic;                                        --  AXI-Stream Receive Data Clk
-----    AXI_STR_RXD_ARESETN     : in  std_logic;                                        --  AXI-Stream Receive Data Reset
-----    AXI_STR_RXD_VALID       : out std_logic;                                        --  AXI-Stream Receive Data Valid
-----    AXI_STR_RXD_READY       : in  std_logic;                                        --  AXI-Stream Receive Data Ready
-----    AXI_STR_RXD_LAST        : out std_logic;                                        --  AXI-Stream Receive Data Last
-----    AXI_STR_RXD_KEEP        : out std_logic_vector(3 downto 0);                     --  AXI-Stream Receive Data Keep
-----    AXI_STR_RXD_DATA        : out std_logic_vector(31 downto 0);                    --  AXI-Stream Receive Data Data
-----
-----    AXI_STR_RXS_ACLK        : in  std_logic;                                        --  AXI-Stream Receive Status Clk
-----    AXI_STR_RXS_ARESETN     : in  std_logic;                                        --  AXI-Stream Receive Status Reset
-----    AXI_STR_RXS_VALID       : out std_logic;                                        --  AXI-Stream Receive Status Valid
-----    AXI_STR_RXS_READY       : in  std_logic;                                        --  AXI-Stream Receive Status Ready
-----    AXI_STR_RXS_LAST        : out std_logic;                                        --  AXI-Stream Receive Status Last
-----    AXI_STR_RXS_KEEP        : out std_logic_vector(3 downto 0);                     --  AXI-Stream Receive Status Keep
-----    AXI_STR_RXS_DATA        : out std_logic_vector(31 downto 0);                    --  AXI-Stream Receive Status Data
-----
-----    -- TEMAC Interface
-----    ------------------------
-----    pause_req               : out std_logic;                                        -- pause req from register to TEMAC
-----    pause_val               : out std_logic_vector(16 to 31);                       -- pause value from register to TEMAC
-----
-----    -- added 05/5/2011
-----    RX_CLK_ENABLE_IN        : in std_logic;                                         -- TEMAC clock domain enable
-----
-----    rx_statistics_vector    : in  std_logic_vector(27 downto 0);                    -- RX statistics from TEMAC
-----    rx_statistics_valid     : in  std_logic;                                        -- Rx stats valid from TEMAC
-----
-----    rx_mac_aclk             : in  std_logic;                                        -- Rx axistream clock from TEMAC
-----    rx_reset                : in  std_logic;                                        -- Rx axistream reset from TEMAC
-----    rx_axis_mac_tdata       : in  std_logic_vector(7 downto 0);                     -- Rx axistream data from TEMAC
-----    rx_axis_mac_tvalid      : in  std_logic;                                        -- Rx axistream valid from TEMAC
-----    rx_axis_mac_tlast       : in  std_logic;                                        -- Rx axistream last from TEMAC
-----    rx_axis_mac_tuser       : in  std_logic;                                        -- Rx axistream good/bad indicator from TEMAC
-----
-----    tx_ifg_delay            : out std_logic_vector(24 to 31);                       -- interframe gap delay from register to TEMAC
-----
-----    tx_mac_aclk             : in  std_logic;                                        -- Tx axistream clock from TEMAC
-----    tx_reset                : in  std_logic;                                        -- Tx axistream reset from TEMAC
-----    tx_axis_mac_tdata       : out std_logic_vector(7 downto 0);                     -- Tx axistream data to TEMAC
-----    tx_axis_mac_tvalid      : out std_logic;                                        -- Tx axistream valid to TEMAC
-----    tx_axis_mac_tlast       : out std_logic;                                        -- Tx axistream last to TEMAC
-----    tx_axis_mac_tuser       : out std_logic;                                        -- Tx axistream underrun indicator to TEMAC
-----    tx_axis_mac_tready      : in  std_logic;                                        -- Tx axistream ready from TEMAC
-----
-----    speed_is_10_100         : in  std_logic;                                        -- speed is 10/100 not 1000 indicator
-----
-----    RESET2TEMAC                     : out std_logic;                                --  Reset to TEMAC
-----
-----    -- Ethernet System signals -----------------------------------------------
-----    PHY_RST_N                       : out std_logic;                                --  Reset to PHY
-----
-----    -- GTX_CLK 125 MHz clock
-----    GTX_CLK                         : in  std_logic                                 --  GTX CLK
-----
-----  );
-----  end component;

-----  component axi_lite_ipif
-----      generic (
-----
-----      C_S_AXI_DATA_WIDTH    : integer  range 32 to 32   := 32;
-----      C_S_AXI_ADDR_WIDTH    : integer                   := 32;
-----      C_S_AXI_MIN_SIZE      : std_logic_vector(31 downto 0):= X"000001FF";
-----      C_USE_WSTRB           : integer := 0;
-----      C_DPHASE_TIMEOUT      : integer range 0 to 512 := 8;
-----      C_ARD_ADDR_RANGE_ARRAY: SLV64_ARRAY_TYPE :=  -- not used
-----      (
-----      X"0000_0000_7000_0000", -- IP user0 base address
-----      X"0000_0000_7000_00FF", -- IP user0 high address
-----      X"0000_0000_7000_0100", -- IP user1 base address
-----      X"0000_0000_7000_01FF"  -- IP user1 high address
-----  );
-----
-----  C_ARD_NUM_CE_ARRAY    : INTEGER_ARRAY_TYPE := -- not used
-----  (
-----  4,         -- User0 CE Number
-----  12         -- User1 CE Number
-----         );
-----         C_FAMILY              : string  := "virtex6"
-----     );
-----     port (
-----
-----      --System signals
-----              S_AXI_ACLK            : in  std_logic;
-----              S_AXI_ARESETN         : in  std_logic;
-----              S_AXI_AWADDR          : in  std_logic_vector (C_S_AXI_ADDR_WIDTH-1 downto 0);
-----              S_AXI_AWVALID         : in  std_logic;
-----              S_AXI_AWREADY         : out std_logic;
-----              S_AXI_WDATA           : in  std_logic_vector (C_S_AXI_DATA_WIDTH-1 downto 0);
-----              S_AXI_WSTRB           : in  std_logic_vector ((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
-----              S_AXI_WVALID          : in  std_logic;
-----              S_AXI_WREADY          : out std_logic;
-----              S_AXI_BRESP           : out std_logic_vector(1 downto 0);
-----              S_AXI_BVALID          : out std_logic;
-----              S_AXI_BREADY          : in  std_logic;
-----              S_AXI_ARADDR          : in  std_logic_vector (C_S_AXI_ADDR_WIDTH-1 downto 0);
-----              S_AXI_ARVALID         : in  std_logic;
-----              S_AXI_ARREADY         : out std_logic;
-----              S_AXI_RDATA           : out std_logic_vector (C_S_AXI_DATA_WIDTH-1 downto 0);
-----              S_AXI_RRESP           : out std_logic_vector(1 downto 0);
-----              S_AXI_RVALID          : out std_logic;
-----              S_AXI_RREADY          : in  std_logic;
-----      -- Controls to the IP/IPIF modules
-----              Bus2IP_Clk            : out std_logic;
-----              Bus2IP_Resetn         : out std_logic;
-----              Bus2IP_Addr           : out std_logic_vector ((C_S_AXI_ADDR_WIDTH-1) downto 0);
-----              Bus2IP_RNW            : out std_logic;
-----              Bus2IP_BE             : out std_logic_vector (((C_S_AXI_DATA_WIDTH/8)-1) downto 0);
-----              Bus2IP_CS             : out std_logic_vector (((C_ARD_ADDR_RANGE_ARRAY'LENGTH)/2-1) downto 0);
-----              Bus2IP_RdCE           : out std_logic_vector ((calc_num_ce(C_ARD_NUM_CE_ARRAY)-1) downto 0);
-----              Bus2IP_WrCE           : out std_logic_vector ((calc_num_ce(C_ARD_NUM_CE_ARRAY)-1) downto 0);
-----              Bus2IP_Data           : out std_logic_vector ((C_S_AXI_DATA_WIDTH-1) downto 0);
-----              IP2Bus_Data           : in  std_logic_vector ((C_S_AXI_DATA_WIDTH-1) downto 0);
-----              IP2Bus_WrAck          : in  std_logic;
-----              IP2Bus_RdAck          : in  std_logic;
-----              IP2Bus_Error          : in  std_logic
-----          );
-----
-----  end component;

end axi_ethernet_buffer_v2_0_25_pack;


-------------------------------------------------------------------------------
-- axi_ethernet_buffer_v2_0_25.vhd
-- Author     : Xilinx Inc.
-------------------------------------------------------------------------------
--
-- *************************************************************************
--
-- (c) Copyright 1998 - 2011 Xilinx, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER

-- rights to the materials distributed herewith. Except as

-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
--
-- *************************************************************************
--
-------------------------------------------------------------------------------
-- Filename:        axi_ethernet_buffer_v2_0_25.vhd
-- Version:         1.0
-- Description:     top level of axi_ethernet_buffer_v2_0_25
--
-------------------------------------------------------------------------------
-- Author:          MSH & MW
-- History:
--  MBR 20/02/12 - took the code from AXI_ETHERNET to create this as a separate
--                 IPXact core.  The original authors of this code are:
--                 Scott Hurt (MSH) and Michael Welter (MW), 2010.
--                 This top level is adapted from the "embedded_top" entity of
--                 AXI_ETHERNET.  Several ports and generics have been cleaned
--                 up (for example the V6EMAC specific syntax has been removed
--                 since the V6 family (and S6 family) are not supported in
--                 Vivado.  I have also replaced C_PHY_TYPE generic with
--                 C_HAS_SGMII (0 or 1).
-- MBR  01/30/2013 - rewritten with better metastability tolerance
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "clk", "clk_div#", "clk_#x"
--      reset signals:                          "rst", "rst_n"
--      generics:                               "C_*"
--      user defined types:                     "*_TYPE"
--      state machine next state:               "*_ns"
--      state machine current state:            "*_cs"
--      combinatorial signals:                  "*_com"
--      pipelined or register delay signals:    "*_d#"
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce"
--      internal version of output port         "*_i"
--      device pins:                            "*_pin"
--      ports:                                  - Names begin with Uppercase
--      processes:                              "*_PROCESS"
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

library axi_lite_ipif_v3_0_5;
use axi_lite_ipif_v3_0_5.all;
use axi_lite_ipif_v3_0_5.ipif_pkg.SLV64_ARRAY_TYPE;
use axi_lite_ipif_v3_0_5.ipif_pkg.INTEGER_ARRAY_TYPE;

library work;
use work.rx_if_pack.all;
use work.tx_if_pack.all;
use work.registers_pack.all;
use work.clock_cross_pack.all;
use work.axi_ethernet_buffer_v2_0_25_pack.all;

-------------------------------------------------------------------------------
-- Definition of Generics :
-------------------------------------------------------------------------------
-- Ethernet generics ??? only requried at the app core level
--  C_TYPE
--     0  Soft TEMAC capable of 10 or 100 Mbps
--     1  Soft TEMAC capable of 10, 100, or 1000 Mbps
--     2  V6 hard TEMAC capable of 10, 100, or 1000 Mbps
--  C_PHY_TYPE
--     0  MII
--     1  GMII
--     2  RGMII V1.3
--     3  RGMII V2.0
--     4  SGMII
--     5  1000Base-X PCS/PMA @ 1 Gbps
--     6  1000Base-X PCS/PMA @ 2 Gbps (C_TYPE=2 only)
--     7  1000Base-X PCS/PMA @ 2.5 Gbps (C_TYPE=2 only)
-------------------------------------------------------------------------------
-- Definition of Generics :
-------------------------------------------------------------------------------
-- System generics
--  C_FAMILY              -- Xilinx FPGA Family
-- AXI generics
--  C_S_AXI_ADDR_WIDTH     -- Width of AXI Address Bus (in bits) 32
--  C_S_AXI_DATA_WIDTH     -- Width of the AXI Data Bus (in bits) 32
--
--  C_HALFDUP             -- Enable half duplex
--  C_TXMEM               -- Depth of TX memory in Bytes
--  C_RXMEM               -- Depth of RX memory in Bytes
--  C_TXCSUM
--     0  No checksum offloading
--     1  Partial (legacy) checksum offloading
--     2  Full checksum offloading
--  C_RXCSUM
--     0  No checksum offloading
--     1  Partial (legacy) checksum offloading
--     2  Full checksum offloading
--  C_TXVLAN_TRAN         -- Enable TX enhanced VLAN translation
--  C_RXVLAN_TRAN         -- Enable RX enhanced VLAN translation
--  C_TXVLAN_TAG          -- Enable TX enhanced VLAN taging
--  C_RXVLAN_TAG          -- Enable RX enhanced VLAN taging
--  C_TXVLAN_STRP         -- Enable TX enhanced VLAN striping
--  C_RXVLAN_STRP         -- Enable RX enhanced VLAN striping
--  C_MCAST_EXTEND        -- Enable RX extended multicast address filtering

-------------------------------------------------------------------------------
--                  Entity Section
-------------------------------------------------------------------------------

entity axi_ethernet_buffer_v2_0_25 is
  generic (
    --  System Generics
    C_FAMILY               : string                        := "virtex7";
    C_S_AXI_ADDR_WIDTH     : integer range 32 to 32        := 32;
    C_S_AXI_DATA_WIDTH     : integer range 32 to 32        := 32;
    C_TEMAC_ADDR_WIDTH     : integer range 0 to 32        := 12;
    C_HALFDUP              : integer range 0 to 1          := 0;
    C_TXMEM                : integer                       := 4096;
    C_RXMEM                : integer                       := 4096;
    C_TXCSUM               : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_RXCSUM               : integer range 0 to 2          := 0;
      -- 0 - No checksum offloading
      -- 1 - Partial (legacy) checksum offloading
      -- 2 - Full checksum offloading
    C_TXVLAN_TRAN          : integer range 0 to 1          := 0;
    C_RXVLAN_TRAN          : integer range 0 to 1          := 0;
    C_TXVLAN_TAG           : integer range 0 to 1          := 0;
    C_RXVLAN_TAG           : integer range 0 to 1          := 0;
    C_TXVLAN_STRP          : integer range 0 to 1          := 0;
    C_RXVLAN_STRP          : integer range 0 to 1          := 0;
    C_MCAST_EXTEND         : integer range 0 to 1          := 0;
    C_SIMULATION           : integer                       := 0;

    C_AVB                 : integer range 0 to 1          := 0;
    C_STATS               : integer range 0 to 1          := 0;
    C_ENABLE_LVDS         : integer range 0 to 1          := 0;
    C_PHY_TYPE            : integer range 0 to 5          := 1;
    C_SPEED_2P5           : integer range 0 to 1          := 0;
    C_PHYADDR             : integer range 0 to 31    := 1; 
    C_PHY_RST_COUNT       : integer   := 1321; 
    C_ENABLE_1588         : integer     := 0;
    C_TYPE                : integer range 0 to 2          := 0
  );
  port (
    -- System signals ---------------------------------------------------------
    S_AXI_ACLK              : in  std_logic;
    S_AXI_ARESETN           : in  std_logic;
    INTERRUPT               : out std_logic;                                        --  AXI Ethernet Interrupt
    -- AXI Lite signals
    S_AXI_AWADDR            : in  std_logic_vector (17 downto 0);
    S_AXI_AWVALID           : in  std_logic;
    S_AXI_AWREADY           : out std_logic;
    S_AXI_WDATA             : in  std_logic_vector  (31 downto 0);
    S_AXI_WSTRB             : in  std_logic_vector (3 downto 0);
    S_AXI_WVALID            : in  std_logic;
    S_AXI_WREADY            : out std_logic;
    S_AXI_BRESP             : out std_logic_vector(1 downto 0);
    S_AXI_BVALID            : out std_logic;
    S_AXI_BREADY            : in  std_logic;
    S_AXI_ARADDR            : in  std_logic_vector (17 downto 0);
    S_AXI_ARVALID           : in  std_logic;
    S_AXI_ARREADY           : out std_logic;
    S_AXI_RDATA             : out std_logic_vector (31 downto 0);
    S_AXI_RRESP             : out std_logic_vector(1 downto 0);
    S_AXI_RVALID            : out std_logic;
    S_AXI_RREADY            : in  std_logic;


    -- Interrupt sources
    EMAC_CLIENT_AUTONEG_INT : in  std_logic;                                        --  Auto negotiation signal from EMAC
    EMAC_RESET_DONE_INT     : in  std_logic;                                        --  Reset Done signal from EMAC
    EMAC_RX_DCM_LOCKED_INT  : in  std_logic;                                        --  DCM Locked signal from EMAC
    PCSPMA_STATUS_VECTOR    : in  std_logic_vector(15 downto 0);                    --  Link Status vector from PCS/PMA core
--    TEMAC_IPIC2GHI_INTR     : in  std_logic;                                        --  Interrupt


    -- AXI Stream signals
    AXI_STR_TXD_ACLK      : in  std_logic;                                          --  AXI-Stream Transmit Data Clk
    AXI_STR_TXD_ARESETN   : in  std_logic;                                          --  AXI-Stream Transmit Data Reset
    AXI_STR_TXD_TVALID    : in  std_logic;                                          --  AXI-Stream Transmit Data Valid
    AXI_STR_TXD_TREADY    : out std_logic;                                          --  AXI-Stream Transmit Data Ready
    AXI_STR_TXD_TLAST     : in  std_logic;                                          --  AXI-Stream Transmit Data Last
    AXI_STR_TXD_TKEEP     : in  std_logic_vector(3 downto 0);                       --  AXI-Stream Transmit Data Keep
    AXI_STR_TXD_TDATA     : in  std_logic_vector(31 downto 0);                      --  AXI-Stream Transmit Data Data

    AXI_STR_TXC_ACLK      : in  std_logic;                                          --  AXI-Stream Transmit Control Clk
    AXI_STR_TXC_ARESETN   : in  std_logic;                                          --  AXI-Stream Transmit Control Reset
    AXI_STR_TXC_TVALID    : in  std_logic;                                          --  AXI-Stream Transmit Control Valid
    AXI_STR_TXC_TREADY    : out std_logic;                                          --  AXI-Stream Transmit Control Ready
    AXI_STR_TXC_TLAST     : in  std_logic;                                          --  AXI-Stream Transmit Control Last
    AXI_STR_TXC_TKEEP     : in  std_logic_vector(3 downto 0);                       --  AXI-Stream Transmit Control Keep
    AXI_STR_TXC_TDATA     : in  std_logic_vector(31 downto 0);                      --  AXI-Stream Transmit Control Data

    AXI_STR_RXD_ACLK        : in  std_logic;                                        --  AXI-Stream Receive Data Clk
    AXI_STR_RXD_ARESETN     : in  std_logic;                                        --  AXI-Stream Receive Data Reset
    AXI_STR_RXD_VALID       : out std_logic;                                        --  AXI-Stream Receive Data Valid
    AXI_STR_RXD_READY       : in  std_logic;                                        --  AXI-Stream Receive Data Ready
    AXI_STR_RXD_LAST        : out std_logic;                                        --  AXI-Stream Receive Data Last
    AXI_STR_RXD_KEEP        : out std_logic_vector(3 downto 0);                     --  AXI-Stream Receive Data Keep
    AXI_STR_RXD_DATA        : out std_logic_vector(31 downto 0);                    --  AXI-Stream Receive Data Data

    AXI_STR_RXS_ACLK        : in  std_logic;                                        --  AXI-Stream Receive Status Clk
    AXI_STR_RXS_ARESETN     : in  std_logic;                                        --  AXI-Stream Receive Status Reset
    AXI_STR_RXS_VALID       : out std_logic;                                        --  AXI-Stream Receive Status Valid
    AXI_STR_RXS_READY       : in  std_logic;                                        --  AXI-Stream Receive Status Ready
    AXI_STR_RXS_LAST        : out std_logic;                                        --  AXI-Stream Receive Status Last
    AXI_STR_RXS_KEEP        : out std_logic_vector(3 downto 0);                     --  AXI-Stream Receive Status Keep
    AXI_STR_RXS_DATA        : out std_logic_vector(31 downto 0);                    --  AXI-Stream Receive Status Data

    -- TEMAC Interface
    ------------------------
    pause_req               : out std_logic;                                        -- pause req from register to TEMAC
    pause_val               : out std_logic_vector(16 to 31);                       -- pause value from register to TEMAC

  ------------------------------
    -- Signals added for axi lite split logic
    S_AXI_2TEMAC_AWADDR : out STD_LOGIC_VECTOR ( C_TEMAC_ADDR_WIDTH - 1 downto 0 );
    S_AXI_2TEMAC_AWVALID : out STD_LOGIC;
    S_AXI_2TEMAC_AWREADY : in STD_LOGIC;
    S_AXI_2TEMAC_WDATA : out STD_LOGIC_VECTOR ( 31 downto 0 );
    S_AXI_2TEMAC_WVALID : out STD_LOGIC;
    S_AXI_2TEMAC_WREADY : in STD_LOGIC;
    S_AXI_2TEMAC_BRESP : in STD_LOGIC_VECTOR ( 1 downto 0 );
    S_AXI_2TEMAC_BVALID : in STD_LOGIC;
    S_AXI_2TEMAC_BREADY : out STD_LOGIC;
    S_AXI_2TEMAC_ARADDR : out STD_LOGIC_VECTOR ( C_TEMAC_ADDR_WIDTH - 1 downto 0 );
    S_AXI_2TEMAC_ARVALID : out STD_LOGIC;
    S_AXI_2TEMAC_ARREADY : in STD_LOGIC;
    S_AXI_2TEMAC_RDATA : in STD_LOGIC_VECTOR ( 31 downto 0 );
    S_AXI_2TEMAC_RRESP : in STD_LOGIC_VECTOR ( 1 downto 0 );
    S_AXI_2TEMAC_RVALID : in STD_LOGIC;
    S_AXI_2TEMAC_RREADY : out STD_LOGIC;
    -- end of Signals added for axi lite split logic
  ------------------------------

    -- added 05/5/2011
    RX_CLK_ENABLE_IN        : in std_logic;                                         -- TEMAC clock domain enable

    rx_statistics_vector    : in  std_logic_vector(27 downto 0);                    -- RX statistics from TEMAC
    rx_statistics_valid     : in  std_logic;                                        -- Rx stats valid from TEMAC

    rx_mac_aclk             : in  std_logic;                                        -- Rx axistream clock from TEMAC
    rx_reset                : in  std_logic;                                        -- Rx axistream reset from TEMAC
    rx_axis_mac_tdata       : in  std_logic_vector(7 downto 0);                     -- Rx axistream data from TEMAC
    rx_axis_mac_tvalid      : in  std_logic;                                        -- Rx axistream valid from TEMAC
    rx_axis_mac_tlast       : in  std_logic;                                        -- Rx axistream last from TEMAC
    rx_axis_mac_tuser       : in  std_logic;                                        -- Rx axistream good/bad indicator from TEMAC

    tx_ifg_delay            : out std_logic_vector(24 to 31);                       -- interframe gap delay from register to TEMAC

    tx_mac_aclk             : in  std_logic;                                        -- Tx axistream clock from TEMAC
    tx_reset                : in  std_logic;                                        -- Tx axistream reset from TEMAC
    tx_axis_mac_tdata       : out std_logic_vector(7 downto 0);                     -- Tx axistream data to TEMAC
    tx_axis_mac_tvalid      : out std_logic;                                        -- Tx axistream valid to TEMAC
    tx_axis_mac_tlast       : out std_logic;                                        -- Tx axistream last to TEMAC
    tx_axis_mac_tuser       : out std_logic_vector(0 downto 0);                                        -- Tx axistream underrun indicator to TEMAC
    tx_axis_mac_tready      : in  std_logic;                                        -- Tx axistream ready from TEMAC
--    tx_collision            : in  std_logic;                                        -- Tx collision not used from TEMAC
--    tx_retransmit           : in  std_logic;                                        -- Tx retransmit not used from TEMAC

    speed_is_10_100         : in  std_logic;                                        -- speed is 10/100 not 1000 indicator

    RESET2PCSPMA                    : out std_logic;                                --  Reset to TEMAC
    RESET2TEMACn                    : out std_logic;                                --  Reset to TEMAC (active low version)

    -- Ethernet System signals -----------------------------------------------
    PHY_RST_N                       : out std_logic;                                --  Reset to PHY

    mdio_i_top    : in   std_logic; -- input from top
    mdio_o_top    : out  std_logic;
    mdio_t_top    : out  std_logic;
    mdc_top       : out  std_logic;
    mdio_t_pcspma : in   std_logic; -- input from pcspma
    mdio_o_pcspma : in   std_logic; -- input from pcspma
    mdio_i_temac  : out  std_logic; -- output to temac
    mdio_o_temac  : in   std_logic;
    mdio_t_temac  : in   std_logic;
    mdc_temac     : in   std_logic;

    -- GTX_CLK 125 MHz clock
    GTX_CLK                         : in  std_logic                                 --  GTX CLK


  );

end axi_ethernet_buffer_v2_0_25;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture imp of axi_ethernet_buffer_v2_0_25 is

    attribute DowngradeIPIdentifiedWarnings: string;
    attribute DowngradeIPIdentifiedWarnings of imp : architecture is "yes";

  ----------------------------------------------------------------------------
  --  Function Declarations
  ----------------------------------------------------------------------------

  function SetVLANWidth (inputTrans, inputStrip, inputTag : integer) return integer is
  Variable vlanWidth : Integer := 1;

    begin
      if (inputTrans = 0 and inputStrip = 0 and inputTag = 0) then
      --  force to be one for lint where in registers.vhd
      --    axiClkTxVlanRdData_i : std_logic_vector(((31-C_TXVLAN_WIDTH)+1) to 31)
      --    bus width would be 32 to 31
        vlanWidth := 1;
      else

        vlanWidth := ((inputTrans*12) + inputStrip + inputTag);
      end if;
    return(vlanWidth);
  end function SetVLANWidth;

  function Set_C_HAS_SGMII (c_phy_type : integer) return integer is
      variable out_val : integer := 0;
    begin
      if (c_phy_type = 4) then
          out_val := 1;
      else
          out_val := 0;
      end if ; 
      return (out_val);
  end function ; 

  ---------------------------------------------------------------------------
  --  Constant Declarations
  ---------------------------------------------------------------------------
  constant C_NUM_CS              : integer := 10;
  constant C_NUM_CE              : integer := 41;
  constant C_SOFT_SIMULATION     : boolean := (C_SIMULATION = 1);
  constant C_TXVLAN_WIDTH : integer := SetVLANWidth(C_TXVLAN_TRAN,C_TXVLAN_STRP,C_TXVLAN_TAG);
  constant C_RXVLAN_WIDTH : integer := SetVLANWidth(C_RXVLAN_TRAN,C_RXVLAN_STRP,C_RXVLAN_TAG);
  --  constant C_TXVLAN_WIDTH : integer := (C_TXVLAN_TRAN*12) + C_TXVLAN_TAG + C_TXVLAN_STRP;
  --  constant C_RXVLAN_WIDTH : integer := (C_RXVLAN_TRAN*12) + C_RXVLAN_TAG + C_RXVLAN_STRP;

    constant C_HAS_SGMII            : integer range 0 to 1          := Set_C_HAS_SGMII(C_PHY_TYPE);

  constant C_ARD_ADDR_RANGE_ARRAY  : SLV64_ARRAY_TYPE :=
    -- Base address and high address pairs.
    (
--      X"00000000" & (C_BASEADDR), -- user0 base address soft registers
--      X"00000000" & (C_HIGHADDR)  -- user0 high address
      X"0000000000000000", -- user0 base address soft registers
      X"000000000003FFFF"  -- user0 high address
    );

  constant C_ARD_NUM_CE_ARRAY   : INTEGER_ARRAY_TYPE :=
    -- This array spcifies the number of Chip Enables (CE) that is
    -- required by the cooresponding baseaddr pair.
    (
      0 =>1
    );

  constant C_S_AXI_MIN_SIZE       : std_logic_vector(31 downto 0) := X"0003FFFF";

  constant C_USE_WSTRB            : integer := 0;

  constant C_DPHASE_TIMEOUT       : integer := 42;

  ---------------------------------------------------------------------------
  -- Signal declarations
  ---------------------------------------------------------------------------
  signal bus2ip_clk_i                 : std_logic;
  signal bus2ip_reset_i               : std_logic;
  signal bus2ip_reset_n_i             : std_logic;

  signal bus2shim_cs                  : std_logic_vector(0 to 0);
  signal bus2shim_rd_ce               : std_logic_vector(0 to 0);
  signal bus2shim_wr_ce               : std_logic_vector(0 to 0);
  signal bus2shim_addr                : std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );
  signal bus2shim_data                : std_logic_vector(0 to C_S_AXI_DATA_WIDTH - 1 );
  signal bus2shim_r_nw                : std_logic;
  signal shim2bus_data                : std_logic_vector (0 to C_S_AXI_DATA_WIDTH - 1 );
  signal shim2bus_wr_ack              : std_logic;
  signal shim2bus_rd_ack              : std_logic;

  signal shim2ip_cs                   : std_logic_vector(0 to C_NUM_CS);
  signal shim2ip_rd_ce                : std_logic_vector(0 to C_NUM_CE);
  signal shim2ip_wr_ce                : std_logic_vector(0 to C_NUM_CE);
  signal shim2ip_addr_i               : std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );
  signal shim2ip_data_i               : std_logic_vector(0 to C_S_AXI_DATA_WIDTH - 1 );
  signal shim2ip_r_nw_i               : std_logic;
  signal ip2shim_data                 : std_logic_vector (0 to C_S_AXI_DATA_WIDTH - 1 );
  signal ip2shim_wr_ack               : std_logic;
  signal ip2shim_rd_ack               : std_logic;
  signal ip2shim_error                : std_logic;

  signal intrpts2reg                  : std_logic_vector(23 to 31);
  signal tx_pause_request             : std_logic;
  signal cr_reg_data                  : std_logic_vector(17 to 31);
  signal tx_pause_reg_data_i          : std_logic_vector(16 to 31);
  signal tx_ifg_delay_i               : std_logic_vector(24 to 31);
  signal is_reg_data                  : std_logic_vector(23 to 31);
  signal ip_reg_data                  : std_logic_vector(23 to 31);
  signal ie_reg_data                  : std_logic_vector(23 to 31);
  signal ttag_reg_data                : std_logic_vector(0 to 31);
  signal rtag_reg_data                : std_logic_vector(0 to 31);
  signal tpid0_reg_data               : std_logic_vector(0 to 31);
  signal tpid1_reg_data               : std_logic_vector(0 to 31);
  signal uawl_reg_data                : std_logic_vector(0 to 31);
  signal uawu_reg_data                : std_logic_vector(16 to 31);
  signal reg_ip2bus_wr_ack            : std_logic;
  signal reg_ip2bus_rd_ack            : std_logic;
  signal reg_ip2bus_data              : std_logic_vector(0 to 31);

  signal reset2axi                    : std_logic;
  signal reset2axi_n                  : std_logic;
  signal reset2axi_str_txd            : std_logic;
  signal reset2axi_str_txc            : std_logic;
  signal reset2axi_str_rxd            : std_logic;
  signal reset2axi_str_rxs            : std_logic;
  signal reset2gtx_clk                : std_logic;

  signal phy_reset_cmplte_intr        : std_logic;

  signal rx_cl_clk_rx_tag_reg_data    : std_logic_vector(0 to 31);
  signal rx_cl_clk_tpid0_reg_data     : std_logic_vector(0 to 31);
  signal rx_cl_clk_tpid1_reg_data     : std_logic_vector(0 to 31);
  signal rx_cl_clk_uawl_reg_data      : std_logic_vector(0 to 31);
  signal rx_cl_clk_uawu_reg_data      : std_logic_vector(16 to 31);
  signal rx_cl_clk_raf_reg_data       : std_logic_vector(17 to 31);

  signal rx_cl_clk_mcast_addr         : std_logic_vector(0 to 14);
  signal rx_cl_clk_mcast_en           : std_logic;
  signal rx_cl_clk_mcast_rd_data      : std_logic_vector(0 to 0);

  signal rx_cl_clk_vlan_addr          : std_logic_vector(0 to 11);
  signal rx_cl_clk_vlan_rd_data       : std_logic_vector(18 to 31);
  signal rx_cl_clk_vlan_bram_en_a     : std_logic;
  signal axiStrTxDClk_vlan_addr       : std_logic_vector(11 downto 0);
  signal axiStrTxDClk_vlan_rd_data    : std_logic_vector(13 downto 0);
  signal axiStrTxDClk_vlan_bram_en_a  : std_logic;

  signal rx_cl_clk_bad_frame_enbl     : std_logic;
  signal rx_cl_clk_emulti_fltr_enbl   : std_logic;
  signal rx_cl_clk_new_fnc_enbl       : std_logic;
  signal rx_cl_clk_brdcast_rej        : std_logic;
  signal rx_cl_clk_mulcast_rej        : std_logic;
  signal rx_cl_clk_vstrp_mode         : std_logic_vector(0 to 1);
  signal rx_cl_clk_vtag_mode          : std_logic_vector(0 to 1);

  signal reset2rx_client              : std_logic;
  signal reset2tx_client              : std_logic;

  signal rxclclk_frame_received_intrpt     : std_logic;
  signal rxclclk_frame_rejected_intrpt     : std_logic;
  signal rxclclk_buffer_mem_overflow_intrpt: std_logic;
  signal axiclk_frame_received_intrpt     : std_logic;
  signal axiclk_frame_rejected_intrpt     : std_logic;
  signal axiclk_buffer_mem_overflow_intrpt: std_logic;

  --  Tx Clock Crossing Signals
  signal tx_cr_reg_data                  : std_logic_vector(4 downto 0);
  signal tx_axi_lite_2_txd_strm_raf_data : std_logic_vector(4 downto 0);
  signal TEMAC_IPIC2GHI_INTR_CROSS       : std_logic;
  signal EMAC_CLIENT_AUTONEG_INT_CROSS   : std_logic;
  signal tx_cmplt_cross                  : std_logic;
  signal EMAC_RX_DCM_LOCKED_CROSS        : std_logic;
  signal EMAC_RESET_DONE_CROSS           : std_logic;
  signal phy_reset_cmplte_intr_cross     : std_logic;
  signal tx_cmplt                        : std_logic;

  signal tpid0_reg_data_cross            : std_logic_vector(15 downto 0);
  signal tpid1_reg_data_cross            : std_logic_vector(15 downto 0);
  signal tpid2_reg_data_cross            : std_logic_vector(15 downto 0);
  signal tpid3_reg_data_cross            : std_logic_vector(15 downto 0);

  signal enable_newFncEn                 : std_logic; --Only perform VLAN when the FLAG = 0xA
  signal cr_reg_data_bit20_sync          : std_logic;
  signal newFncEn_cross                  : std_logic;
  signal transMode_cross                 : std_logic;
  signal tagMode_cross                   : std_logic_vector( 1 downto 0);
  signal strpMode_cross                  : std_logic_vector( 1 downto 0);

  signal tpid0_cross                     : std_logic_vector(15 downto 0);
  signal tpid1_cross                     : std_logic_vector(15 downto 0);
  signal tpid2_cross                     : std_logic_vector(15 downto 0);
  signal tpid3_cross                     : std_logic_vector(15 downto 0);

  signal newTagData_cross                : std_logic_vector(31 downto 0);

  signal pcspma_status_cross             : std_logic_vector(16 to 31);

  signal tx_init_in_prog                 : std_logic;
  signal tx_init_in_prog_cross           : std_logic;

    ------------------------------
    -- Signals added for axi lite split logic
    signal valid_awaddr_range      : std_logic_vector (17 downto 0);
    signal valid_awaddr_init_range : std_logic                     ;
    signal valid_araddr_range      : std_logic_vector (17 downto 0);
    signal embedded_araddr         : std_logic                     ;
    signal embedded_araddr1        : std_logic                     ;
    signal embedded_araddr2        : std_logic                     ;
    signal embedded_araddr3        : std_logic                     ;
    signal embedded_araddr_reg     : std_logic                     ;
    signal embedded_araddr_sel     : std_logic                     ;
    signal embedded_awaddr         : std_logic                     ;
    signal embedded_awaddr1        : std_logic                     ;
    signal embedded_awaddr2        : std_logic                     ;
    signal embedded_awaddr3        : std_logic                     ;
    signal embedded_awaddr_reg     : std_logic                     ;
    signal embedded_awaddr_sel     : std_logic                     ;
    signal S_AXI_2EMBED_WVALID     : std_logic                     ;
    signal S_AXI_2EMBED_AWVALID    : std_logic                     ;
    signal S_AXI_2EMBED_ARVALID    : std_logic                     ;
    signal s_axi_awready_embed     : std_logic                     ;
    signal s_axi_wready_embed      : std_logic                     ;
    signal s_axi_bresp_embed       : std_logic_vector ( 1 downto 0);
    signal s_axi_bvalid_embed      : std_logic                     ;
    signal s_axi_arready_embed     : std_logic                     ;
    signal s_axi_rdata_embed       : std_logic_vector (31 downto 0);
    signal s_axi_rresp_embed       : std_logic_vector ( 1 downto 0);
    signal s_axi_rvalid_embed      : std_logic                     ;

    ------------------------------
    -- 01/30/13: new signals for metastability improvements
	signal bus2ip_reset_reg        : std_logic := '0'              ;
	signal sample_config           : std_logic := '0'              ;
    signal sample_rx_mac_config    : std_logic                     ;
    signal sample_tx_mac_config    : std_logic                     ;
    signal sample_axi_str_config   : std_logic                     ;

    signal s_axi_awaddr_int_sig    : std_logic_vector (31 downto 0);
    signal s_axi_araddr_int_sig    : std_logic_vector (31 downto 0);
    signal mdio_t_passthrough   : std_logic                     ;
    signal mdio_o_passthrough   : std_logic                     ;
    signal mdc_passthrough   : std_logic                     ;

begin

  rx_cl_clk_bad_frame_enbl   <= rx_cl_clk_raf_reg_data(17);
  rx_cl_clk_emulti_fltr_enbl <= rx_cl_clk_raf_reg_data(19);
  rx_cl_clk_new_fnc_enbl     <= rx_cl_clk_raf_reg_data(20);
  rx_cl_clk_vstrp_mode       <= rx_cl_clk_raf_reg_data(21 to 22);
  rx_cl_clk_vtag_mode        <= rx_cl_clk_raf_reg_data(25 to 26);
  rx_cl_clk_brdcast_rej      <= rx_cl_clk_raf_reg_data(29);
  rx_cl_clk_mulcast_rej      <= rx_cl_clk_raf_reg_data(30);


--  intrpts2reg(31) <= TEMAC_IPIC2GHI_INTR_CROSS;
  intrpts2reg(31) <= '0';

  intrpts2reg(30) <= EMAC_CLIENT_AUTONEG_INT_CROSS;
  intrpts2reg(29) <= axiclk_frame_received_intrpt; --rx complete
  intrpts2reg(28) <= axiclk_frame_rejected_intrpt; --rx reject
  intrpts2reg(27) <= axiclk_buffer_mem_overflow_intrpt; --rx mem overflow
  intrpts2reg(26) <= tx_cmplt_cross;    --'0'; --tx_cmplt_cross --fix mee - need to implement!!!!!
  intrpts2reg(25) <= EMAC_RX_DCM_LOCKED_CROSS;
  intrpts2reg(24) <= EMAC_RESET_DONE_CROSS;
  intrpts2reg(23) <= phy_reset_cmplte_intr_cross;

  RXCLCLK2AXICLK_INTRPT0 : actv_hi_pulse_clk_cross
  port map    (
    ClkA               => rx_mac_aclk,
    ClkARst            => reset2rx_client,
    ClkASignalIn       => rxclclk_frame_received_intrpt,
    ClkB               => bus2ip_clk_i,
    ClkBRst            => reset2axi,
    ClkBSignalOut      => axiclk_frame_received_intrpt
  );

  RXCLCLK2AXICLK_INTRPT1 : actv_hi_pulse_clk_cross
  port map    (
    ClkA               => rx_mac_aclk,
    ClkARst            => reset2rx_client,
    ClkASignalIn       => rxclclk_frame_rejected_intrpt,
    ClkB               => bus2ip_clk_i,
    ClkBRst            => reset2axi,
    ClkBSignalOut      => axiclk_frame_rejected_intrpt
  );

  RXCLCLK2AXICLK_INTRPT2 : actv_hi_pulse_clk_cross
  port map    (
    ClkA               => rx_mac_aclk,
    ClkARst            => reset2rx_client,
    ClkASignalIn       => rxclclk_buffer_mem_overflow_intrpt,
    ClkB               => bus2ip_clk_i,
    ClkBRst            => reset2axi,
    ClkBSignalOut      => axiclk_buffer_mem_overflow_intrpt
  );


  COMBINE_RESETS : reset_combiner
  generic map (
    C_PHY_RST_COUNT    => C_PHY_RST_COUNT,
    C_FAMILY           => C_FAMILY,
    C_SIMULATION       => C_SIMULATION
  )
  port map    (
    S_AXI_ACLK           => S_AXI_ACLK,
    S_AXI_ARESETN        => S_AXI_ARESETN,
    GTX_CLK_125MHZ       => GTX_CLK,
    RX_CLIENT_CLK        => rx_mac_aclk,
    RX_CLIENT_CLK_EN     => '1', --RX_CLIENT_CLK_ENBL,
    TX_CLIENT_CLK        => tx_mac_aclk,
    TX_CLIENT_CLK_EN     => '1', --TX_CLIENT_CLK_ENBL,
    AXI_STR_TXD_ACLK     => AXI_STR_TXD_ACLK,
    AXI_STR_TXD_ARESETN  => AXI_STR_TXD_ARESETN,
    AXI_STR_TXC_ACLK     => AXI_STR_TXC_ACLK,
    AXI_STR_TXC_ARESETN  => AXI_STR_TXC_ARESETN,
    AXI_STR_RXD_ACLK     => AXI_STR_RXD_ACLK,
    AXI_STR_RXD_ARESETN  => AXI_STR_RXD_ARESETN,
    AXI_STR_RXS_ACLK     => AXI_STR_RXS_ACLK,
    AXI_STR_RXS_ARESETN  => AXI_STR_RXS_ARESETN,
    PHY_RESET_N          => PHY_RST_N, -- >= 10mS as req'd by PHY spec
    PHY_RESET_CMPLTE     => phy_reset_cmplte_intr, -- >= 15mS as req'd by PHY spec
    RESET2AXI            => reset2axi,
    RESET2RX_CLIENT      => reset2rx_client,
    RESET2TX_CLIENT      => reset2tx_client,
    RESET2AXI_STR_TXD    => reset2axi_str_txd,
    RESET2AXI_STR_TXC    => reset2axi_str_txc,
    RESET2AXI_STR_RXD    => reset2axi_str_rxd,
    RESET2AXI_STR_RXS    => reset2axi_str_rxs,
    reset2gtx_clk        => reset2gtx_clk
  );

  reset2axi_n      <= not(reset2axi);
--  RESET2STATISTICS <= reset2axi;
  RESET2PCSPMA      <= reset2axi;
  RESET2TEMACn     <= not reset2axi;
  --------------------------------------------------------------------------
  -- REG_RD_WR_DATA_PROCESS
  --------------------------------------------------------------------------
  REG_RD_WR_DATA_PROCESS : process (bus2ip_clk_i)
  begin
    if (bus2ip_clk_i'event and bus2ip_clk_i = '1') then
      if (bus2ip_reset_i = '1') then
        ip2shim_data   <= (others => '0');
        ip2shim_rd_ack <= '0';
        ip2shim_wr_ack <= '0';
      else
        ip2shim_data   <= reg_ip2bus_data;
        ip2shim_rd_ack <= reg_ip2bus_rd_ack;
        ip2shim_wr_ack <= reg_ip2bus_wr_ack;

      end if;
    end if;
  end process;
  ip2shim_error  <= '0';


  I_REGISTERS : registers
  generic map (
    C_FAMILY       => C_FAMILY,
    C_TXVLAN_TRAN  => C_TXVLAN_TRAN,
    C_TXVLAN_TAG   => C_TXVLAN_TAG,
    C_TXVLAN_STRP  => C_TXVLAN_STRP,
    C_RXVLAN_TRAN  => C_RXVLAN_TRAN,
    C_RXVLAN_TAG   => C_RXVLAN_TAG,
    C_RXVLAN_STRP  => C_RXVLAN_STRP,
    C_MCAST_EXTEND => C_MCAST_EXTEND,
    C_TXVLAN_WIDTH => C_TXVLAN_WIDTH,
    C_RXVLAN_WIDTH => C_RXVLAN_WIDTH
  )
  port map    (
    AxiClk                    => bus2ip_clk_i,      -- in
    AXI_STR_TXD_ACLK          => AXI_STR_TXD_ACLK,
    RxClClk                   => rx_mac_aclk,   --: in
    AxiReset                  => bus2ip_reset_i,     -- in  from top level system
    IP2BUS_DATA               => reg_ip2bus_data, -- out to shim
    IP2Bus_WrAck              => reg_ip2bus_wr_ack,-- out to shim
    IP2Bus_RdAck              => reg_ip2bus_rd_ack,-- out to shim
    BUS2IP_ADDR               => shim2ip_addr_i,    -- in  from shim
    BUS2IP_DATA               => shim2ip_data_i,    -- in  from shim
    Bus2IP_RNW                => shim2ip_r_nw_i,    -- in  from shim
    BUS2IP_CS                 => shim2ip_cs  ,    -- in  from shim
    Bus2IP_RdCE               => shim2ip_rd_ce,    -- in  from shim
    Bus2IP_WrCE               => shim2ip_wr_ce,    -- in  from shim
    IntrptsIn                 => intrpts2reg,    -- in
    TPReq                     => tx_pause_request,           -- out
    CrRegData                 => cr_reg_data,       -- out
    TpRegData                 => tx_pause_reg_data_i,       -- out
    IfgpRegData               => tx_ifg_delay_i,     -- out
    IsRegData                 => is_reg_data,       -- out
    IpRegData                 => ip_reg_data,       -- out
    IeRegData                 => ie_reg_data,       -- out
    IntrptOut                 => INTERRUPT,       -- out
    TtagRegData               => ttag_reg_data,     -- out
    RtagRegData               => rtag_reg_data,     -- out
    Tpid0RegData              => tpid0_reg_data,    -- out
    Tpid1RegData              => tpid1_reg_data,    -- out
    pcspma_status_cross       => pcspma_status_cross,
    UawLRegData               => uawl_reg_data,           -- out
    UawURegData               => uawu_reg_data,           -- out
    RxClClkMcastAddr          => rx_cl_clk_mcast_addr,      -- in
    RxClClkMcastEn            => rx_cl_clk_mcast_en,        -- in
    RxClClkMcastRdData        => rx_cl_clk_mcast_rd_data,    -- out
    AxiStrTxDClkTxVlanAddr    => axiStrTxDClk_vlan_addr,   -- in
    AxiStrTxDClkTxVlanRdData  => axiStrTxDClk_vlan_rd_data, -- out
    RxClClkRxVlanAddr         => rx_cl_clk_vlan_addr,   -- in
    RxClClkRXVlanRdData       => rx_cl_clk_vlan_rd_data, -- out
    AxiStrTxDClkTxVlanBramEnA => axiStrTxDClk_vlan_bram_en_a,-- in
    RxClClkRxVlanBramEnA      => rx_cl_clk_vlan_bram_en_a -- in
  );


    ------------------------------
    -- Logic added for axi lite split functionality

    valid_araddr_range <= S_AXI_ARADDR (17 downto 0);
    embedded_araddr_sel <=  embedded_araddr when (S_AXI_ARVALID = '1') else embedded_araddr_reg ;
    embedded_araddr <=  embedded_araddr1 OR embedded_araddr2 OR embedded_araddr3;
    embedded_araddr1 <=  '1' when (valid_araddr_range >= "000000000000000000" and valid_araddr_range <= "000000000000110000" ) else '0';
    embedded_araddr2 <=  '1' when (valid_araddr_range(17 downto 14) = "0001" or valid_araddr_range(17 downto 14) = "0010" ) else '0';
    embedded_araddr3 <=  '1' when (valid_araddr_range(17) = '1') else '0';
    embedded_araddr_reg_process : process (S_AXI_ACLK)
    begin
      if (S_AXI_ACLK'event and S_AXI_ACLK = '1') then
          if (S_AXI_ARESETN = '0') then
              embedded_araddr_reg    <= '0';
          else
              embedded_araddr_reg    <= embedded_araddr_sel;
          end if;
      end if;
    end process;

    valid_awaddr_range <= S_AXI_AWADDR (17 downto 0);
    embedded_awaddr_sel <=  embedded_awaddr when (S_AXI_AWVALID = '1') else embedded_awaddr_reg ;
    embedded_awaddr <=  embedded_awaddr1 OR embedded_awaddr2 OR embedded_awaddr3;
    embedded_awaddr1 <=  '1' when (valid_awaddr_range >= "000000000000000000" and valid_awaddr_range <= "000000000000110000" ) else '0';
    embedded_awaddr2 <=  '1' when (valid_awaddr_range(17 downto 14) = "0001" or valid_awaddr_range(17 downto 14) = "0010" ) else '0';
    embedded_awaddr3 <=  '1' when (valid_awaddr_range(17) = '1') else '0';
    embedded_awaddr_reg_process : process (S_AXI_ACLK)
    begin
      if (S_AXI_ACLK'event and S_AXI_ACLK = '1') then
          if (S_AXI_ARESETN = '0') then
              embedded_awaddr_reg    <= '0';
          else
              embedded_awaddr_reg    <= embedded_awaddr_sel;
          end if;
      end if;
    end process;

    S_AXI_2TEMAC_AWADDR  <= s_axi_awaddr(C_TEMAC_ADDR_WIDTH -1  downto 0); 
    S_AXI_2TEMAC_AWVALID <= s_axi_awvalid and not embedded_awaddr_sel; -- : out STD_LOGIC;
    S_AXI_2TEMAC_WDATA   <= s_axi_wdata; -- : out STD_LOGIC_VECTOR ( 31 downto 0 );
    S_AXI_2TEMAC_WVALID  <= s_axi_wvalid and not embedded_awaddr_sel; -- : out STD_LOGIC;
    S_AXI_2TEMAC_BREADY  <= s_axi_bready; -- : out STD_LOGIC;
    S_AXI_2TEMAC_ARADDR  <= s_axi_araddr(C_TEMAC_ADDR_WIDTH -1  downto 0);
    S_AXI_2TEMAC_ARVALID <= s_axi_arvalid and not embedded_araddr_sel; -- : out STD_LOGIC;
    S_AXI_2TEMAC_RREADY  <= s_axi_rready; -- : out STD_LOGIC;

    S_AXI_2EMBED_WVALID  <= s_axi_wvalid and embedded_awaddr_sel; -- : out STD_LOGIC;
    S_AXI_2EMBED_AWVALID <= s_axi_awvalid and embedded_awaddr_sel; -- : out STD_LOGIC;
    S_AXI_2EMBED_ARVALID <= s_axi_arvalid and embedded_araddr_sel; -- : out STD_LOGIC;

    s_axi_awready <= s_axi_awready_embed  when ( embedded_awaddr_sel = '1' ) else  S_AXI_2TEMAC_AWREADY ; --: in STD_LOGIC  ;
    s_axi_wready  <= s_axi_wready_embed   when ( embedded_awaddr_sel = '1' ) else  S_AXI_2TEMAC_WREADY  ; --: in STD_LOGIC  ;
    s_axi_bresp   <= s_axi_bresp_embed    when ( embedded_awaddr_sel = '1' ) else  S_AXI_2TEMAC_BRESP   ; --: in STD_LOGIC_VECTOR ( 1 downto 0 )  ;
    s_axi_bvalid  <= s_axi_bvalid_embed   when ( embedded_awaddr_sel = '1' ) else  S_AXI_2TEMAC_BVALID  ; --: in STD_LOGIC  ;
    s_axi_arready <= s_axi_arready_embed  when ( embedded_araddr_sel = '1' ) else  S_AXI_2TEMAC_ARREADY ; --: in STD_LOGIC  ;
    s_axi_rdata   <= s_axi_rdata_embed    when ( embedded_araddr_sel = '1' ) else  S_AXI_2TEMAC_RDATA   ; --: in STD_LOGIC_VECTOR ( 31 downto 0 ) ;
    s_axi_rresp   <= s_axi_rresp_embed    when ( embedded_araddr_sel = '1' ) else  S_AXI_2TEMAC_RRESP   ; --: in STD_LOGIC_VECTOR ( 1 downto 0 )  ;
    s_axi_rvalid  <= s_axi_rvalid_embed   when ( embedded_araddr_sel = '1' ) else  S_AXI_2TEMAC_RVALID  ; --: in STD_LOGIC  ;

  -- End of logic added for axi lite split logic
    ------------------------------

  --------------------------------------------------------------------------
  -- Instantiate AXI lite IPIF
  --------------------------------------------------------------------------
    s_axi_awaddr_int_sig   <=  "00000000000000" & S_AXI_AWADDR;
    s_axi_araddr_int_sig   <=  "00000000000000" & S_AXI_ARADDR;

  I_AXI_LITE_IPIF : entity axi_lite_ipif_v3_0_5.axi_lite_ipif
  generic map (
    C_FAMILY                  => C_FAMILY,
    C_S_AXI_ADDR_WIDTH        => C_S_AXI_ADDR_WIDTH,
    C_S_AXI_DATA_WIDTH        => C_S_AXI_DATA_WIDTH,
    C_S_AXI_MIN_SIZE          => C_S_AXI_MIN_SIZE,
    C_USE_WSTRB               => C_USE_WSTRB,
    C_DPHASE_TIMEOUT          => C_DPHASE_TIMEOUT,
    C_ARD_ADDR_RANGE_ARRAY    => C_ARD_ADDR_RANGE_ARRAY,
    C_ARD_NUM_CE_ARRAY        => C_ARD_NUM_CE_ARRAY
  )
  port map (
    S_AXI_ACLK     =>  S_AXI_ACLK,
    S_AXI_ARESETN  =>  reset2axi_n,
    S_AXI_AWADDR   =>  s_axi_awaddr_int_sig,
    S_AXI_AWVALID  =>  S_AXI_2EMBED_AWVALID,
    S_AXI_AWREADY  =>  S_AXI_AWREADY_embed,
    S_AXI_WDATA    =>  S_AXI_WDATA,
    S_AXI_WSTRB    =>  S_AXI_WSTRB,
    S_AXI_WVALID   =>  S_AXI_2EMBED_WVALID,
    S_AXI_WREADY   =>  S_AXI_WREADY_embed,
    S_AXI_BRESP    =>  S_AXI_BRESP_embed,
    S_AXI_BVALID   =>  S_AXI_BVALID_embed,
    S_AXI_BREADY   =>  S_AXI_BREADY,
    S_AXI_ARADDR   =>  s_axi_araddr_int_sig,
    S_AXI_ARVALID  =>  S_AXI_2EMBED_ARVALID,
    S_AXI_ARREADY  =>  S_AXI_ARREADY_embed,
    S_AXI_RDATA    =>  S_AXI_RDATA_embed,
    S_AXI_RRESP    =>  S_AXI_RRESP_embed,
    S_AXI_RVALID   =>  S_AXI_RVALID_embed,
    S_AXI_RREADY   =>  S_AXI_RREADY,

    -- IP Interconnect (IPIC) port signals
    BUS2IP_CLK     => bus2ip_clk_i,
    BUS2IP_RESETN  => bus2ip_reset_n_i,
    IP2BUS_DATA    => shim2bus_data ,
    IP2BUS_WRACK   => shim2bus_wr_ack,
    IP2BUS_RDACK   => shim2bus_rd_ack,
    IP2BUS_ERROR   => ip2shim_error,
    BUS2IP_ADDR    => bus2shim_addr,
    BUS2IP_DATA    => bus2shim_data,
    BUS2IP_RNW     => bus2shim_r_nw ,
    BUS2IP_BE      => open,
    BUS2IP_CS      => bus2shim_cs  ,
    BUS2IP_RDCE    => bus2shim_rd_ce,
    BUS2IP_WRCE    => bus2shim_wr_ce
  );

 bus2ip_reset_i <= not(bus2ip_reset_n_i);
--  bus2ip_reset_i <= not(reset2axi_n);

  -- Instantiate the Address response shim for invalid addresses
  I_ADDR_SHIM : addr_response_shim
  generic map(
    C_BUS2CORE_CLK_RATIO      => 1,
    C_S_AXI_ADDR_WIDTH        => C_S_AXI_ADDR_WIDTH,
    C_S_AXI_DATA_WIDTH        => C_S_AXI_DATA_WIDTH,
    C_SIPIF_DWIDTH            => 32,
    C_NUM_CS                  => C_NUM_CS,
    C_NUM_CE                  => C_NUM_CE,
    C_FAMILY                  => C_FAMILY
  )
  port map(
    -- clock and reset                                    -- --Clock and Reset
    BUS2IP_CLK                => bus2ip_clk_i,            -- : in  std_logic;                                        --  AXI4-Lite clk
    BUS2IP_RESET              => bus2ip_reset_i,          -- : in  std_logic;                                        --  AXI4-Lite reset
                                                          --
    -- slave AXI bus interface with shim                  -- -- PLB Slave Interface with Shim
    BUS2IP_ADDR             =>  bus2shim_addr, -- BUS2IP_ADDR,               -- : in  std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );   --  Address bus from AXI4-Lite to Shim
    BUS2IP_DATA             =>  bus2shim_data, -- BUS2IP_DATA,               -- : in  std_logic_vector(0 to C_SIPIF_DWIDTH - 1 );       --  Data bus from AXI4-Lite to Shim
    BUS2IP_RNW              =>  bus2shim_r_nw, -- BUS2IP_R_NW ,              -- : in  std_logic;                                        --  RNW signal from AXI4-Lite to Shim
    BUS2IP_CS               =>  bus2shim_cs, -- BUS2IP_CS  ,               -- : in  std_logic_vector(0 to 0);                         --  CS signal from AXI4-Lite to Shim
    BUS2IP_RDCE             =>  bus2shim_rd_ce, -- BUS2IP_RDCE,               -- : in  std_logic_vector(0 to 0);                         --  RdCE signal from AXI4-Lite to Shim
    BUS2IP_WRCE             =>  bus2shim_wr_ce, -- BUS2IP_WRCE,               -- : in  std_logic_vector(0 to 0);                         --  WrCE signal from AXI4-Lite to Shim
                                 --                            --
    IP2BUS_DATA             =>  shim2bus_data, -- IP2BUS_DATA ,              -- : out std_logic_vector (0 to C_SIPIF_DWIDTH - 1 );      --  Data bus from Shim to AXI4-Lite
    IP2BUS_WRACK            =>  shim2bus_wr_ack, -- IP2BUS_WR_ACK,             -- : out std_logic;                                        --  WrCE signal from Shim to AXI4-Lite
    IP2BUS_RDACK            =>  shim2bus_rd_ack, -- IP2BUS_RD_ACK,             -- : out std_logic;                                        --  RdCE signal from Shim to AXI4-Lite
                                                          --
    -- internal interface with shim                       -- -- TEMAC Interface with Shim
    SHIM2IP_ADDR              => shim2ip_addr_i,          -- : out std_logic_vector(0 to C_S_AXI_ADDR_WIDTH - 1 );   --  Address bus from Shim to AXI Ethernet
    SHIM2IP_DATA              => shim2ip_data_i,          -- : out std_logic_vector(0 to C_SIPIF_DWIDTH - 1 );       --  Data bus from Shim to AXI Ethernet
    SHIM2IP_RNW               => shim2ip_r_nw_i,          -- : out std_logic;                                        --  RNW signal from Shim to AXI Ethernet
    SHIM2IP_CS                => shim2ip_cs  ,            -- : out std_logic_vector(0 to C_NUM_CS);                  --  CS signal from Shim to AXI Ethernet
    SHIM2IP_RDCE              => shim2ip_rd_ce,           -- : out std_logic_vector(0 to C_NUM_CE);                  --  RdCE signal from Shim to AXI Ethernet
    SHIM2IP_WRCE              => shim2ip_wr_ce,           -- : out std_logic_vector(0 to C_NUM_CE);                  --  WrCE signal from Shim to AXI Ethernet
                                                          --
    IP2SHIM_DATA              => ip2shim_data,            -- : in  std_logic_vector (0 to C_SIPIF_DWIDTH - 1 );      --  Data bus from AXI Ethernet to Shim
    IP2SHIM_WRACK             => ip2shim_wr_ack,          -- : in  std_logic;                                        --  WrCE signal from AXI Ethernet to Shim
    IP2SHIM_RDACK             => ip2shim_rd_ack           -- : in  std_logic                                         --  RdCE signal from AXI Ethernet to Shim
  );


  -- -------------------------
  -- Here the sample_config signal is created.  This will pulse high after an AXI_Lite clock write
  -- to configuration OR following an AXI-Lite reset (when the configuration is set back to reset
  -- defaults).
  --
  -- The sample_config is then synchronised into an appropriate clock domain to ensure that 
  -- that the configuration data will be stable to sample in the new clock domain.
  -- -------------------------

  gen_sample_config : process (bus2ip_clk_i)
  begin
      if (bus2ip_clk_i'event and bus2ip_clk_i = '1') then
	    bus2ip_reset_reg <= bus2ip_reset_i;
		sample_config    <= reg_ip2bus_wr_ack or (not bus2ip_reset_i and bus2ip_reset_reg);
      end if;
  end process gen_sample_config;

  gen_sample_rx_mac_config : actv_hi_pulse_clk_cross
  port map    (
    ClkA               => bus2ip_clk_i,
    ClkARst            => '0',
    ClkASignalIn       => sample_config,
    ClkB               => rx_mac_aclk,
    ClkBRst            => '0', -- do not use resets here
    ClkBSignalOut      => sample_rx_mac_config
  );

  gen_sample_tx_mac_config : actv_hi_pulse_clk_cross
  port map    (
    ClkA               => bus2ip_clk_i,
    ClkARst            => '0',
    ClkASignalIn       => sample_config,
    ClkB               => tx_mac_aclk,
    ClkBRst            => '0', -- do not use resets here
    ClkBSignalOut      => sample_tx_mac_config
  );

  gen_sample_axi_str_config : actv_hi_pulse_clk_cross
  port map    (
    ClkA               => bus2ip_clk_i,
    ClkARst            => '0',
    ClkASignalIn       => sample_config,
    ClkB               => AXI_STR_TXD_ACLK,
    ClkBRst            => '0', -- do not use resets here
    ClkBSignalOut      => sample_axi_str_config
  );
  -- -------------------------


  TAG_REG_CROSS_I : bus_clk_cross
  generic map (
    C_BUS_WIDTH  => 32
  )
  port map(
    Clk_A_BUS_IN    =>  rtag_reg_data,
    Clk_B           =>  rx_mac_aclk,
    Clk_B_Rst       =>  reset2rx_client,
    stable_for_sample => sample_rx_mac_config,
    ClkBBusOut   =>  rx_cl_clk_rx_tag_reg_data
  );

  TPID0_REG_CROSS_I : bus_clk_cross
  generic map (
    C_BUS_WIDTH  => 32
  )
  port map(
    Clk_A_BUS_IN    =>  tpid0_reg_data,
    Clk_B           =>  rx_mac_aclk,
    Clk_B_Rst       =>  reset2rx_client,
    stable_for_sample => sample_rx_mac_config,
    ClkBBusOut   =>  rx_cl_clk_tpid0_reg_data
  );

  TPID1_REG_CROSS_I : bus_clk_cross
  generic map (
    C_BUS_WIDTH  => 32
  )
  port map(
    Clk_A_BUS_IN    =>  tpid1_reg_data,
    Clk_B           =>  rx_mac_aclk,
    Clk_B_Rst       =>  reset2rx_client,
    stable_for_sample => sample_rx_mac_config,
    ClkBBusOut   =>  rx_cl_clk_tpid1_reg_data
  );

  UAWL_REG_CROSS_I : bus_clk_cross
  generic map (
    C_BUS_WIDTH  => 32
  )
  port map(
    Clk_A_BUS_IN    =>  uawl_reg_data,
    Clk_B           =>  rx_mac_aclk,
    Clk_B_Rst       =>  reset2rx_client,
    stable_for_sample => sample_rx_mac_config,
    ClkBBusOut   =>  rx_cl_clk_uawl_reg_data
  );

  UAWU_REG_CROSS_I : bus_clk_cross
  generic map (
    C_BUS_WIDTH  => 16
  )
  port map(
    Clk_A_BUS_IN    =>  uawu_reg_data,
    Clk_B           =>  rx_mac_aclk,
    Clk_B_Rst       =>  reset2rx_client,
    stable_for_sample => sample_rx_mac_config,
    ClkBBusOut   =>  rx_cl_clk_uawu_reg_data
  );

  RAF_REG_CROSS_I : bus_clk_cross
  generic map (
    C_BUS_WIDTH  => 15
  )
  port map(
    Clk_A_BUS_IN    =>  cr_reg_data,
    Clk_B           =>  rx_mac_aclk,
    Clk_B_Rst       =>  reset2rx_client,
    stable_for_sample => sample_rx_mac_config,
    ClkBBusOut   =>  rx_cl_clk_raf_reg_data
  );

  PCSPMA_STATUS_CROSS_I: for i in 15 downto 0 generate
     sync_pcspma_status: sync_block
     port map (
        clk       => bus2ip_clk_i,
        reset     => reset2axi,
        data_in   => pcspma_status_vector(i),
        data_out  => pcspma_status_cross(31-i)
     );
  end generate;



----------------------------------------------------------------------------
--  Tx Interface Clock Crossing - Start
----------------------------------------------------------------------------

  GEN_TX_VLAN_NEWFNCEN_CROSS : if C_TXVLAN_STRP = 1 or C_TXVLAN_TAG = 1 or C_TXVLAN_TRAN = 1 generate
  begin

    gen_cr_reg_data_bit20_sync : sync_block
    port map (
      clk        => AXI_STR_TXD_ACLK,
      reset      => reset2axi_str_txd,
      data_in    => cr_reg_data(20),
      data_out   => cr_reg_data_bit20_sync
    );

    -- ****** martinr **** check assumption that AXI_STR_TXD_ACLK = AXI_STR_TXC_ACLK
    --  RAF Register Clock crossing
    newFncEn_cross <= cr_reg_data_bit20_sync and enable_newFncEn;          --  NewFncEnbl
  end generate;


  GEN_NO_TX_VLAN_NEWFNCEN_CROSS : if not(C_TXVLAN_STRP = 1 or C_TXVLAN_TAG = 1 or C_TXVLAN_TRAN = 1) generate
  begin

    newFncEn_cross <= '0';
  end generate;


  GEN_TX_VLAN_TRANS_ENABLE : if C_TXVLAN_TRAN = 1 generate
  begin

    transMode_cross <= newFncEn_cross;
  end generate;

  GEN_NO_TX_VLAN_TRANS_ENABLE : if C_TXVLAN_TRAN = 0 generate
  begin

    transMode_cross <= '0';
  end generate;




  GEN_TX_VLAN_STRP_CROSS : if C_TXVLAN_STRP = 1 generate
    signal tx_StripMode : std_logic_vector(1 downto 0);
    signal reset_strp   : std_logic;
  begin

    tx_StripMode  <= cr_reg_data(23 to 24);    --  TxVStripMode
    reset_strp    <= reset2axi_str_txd or not newFncEn_cross;

    TX_STRP_CROSS_I : bus_clk_cross
    generic map (
      C_BUS_WIDTH  => 2
    )
    port map(
      Clk_A_BUS_IN    =>  tx_StripMode,
      Clk_B           =>  AXI_STR_TXD_ACLK,
      Clk_B_Rst       =>  reset_strp,
      stable_for_sample => sample_axi_str_config,
      ClkBBusOut   =>  strpMode_cross
    );
  end generate;

  GEN_NO_TX_VLAN_STRP_CROSS : if C_TXVLAN_STRP = 0 generate
  begin
    strpMode_cross <= (others => '0');
  end generate;


  GEN_TX_VLAN_TAG_CROSS : if C_TXVLAN_TAG = 1 generate
    signal tx_TagMode : std_logic_vector(1 downto 0);
    signal reset_tag  : std_logic;
  begin

    tx_TagMode   <= cr_reg_data(27 to 28);    --  TxVTagMode
    reset_tag    <= reset2axi_str_txd or not newFncEn_cross;

    TX_STRP_CROSS_I : bus_clk_cross
    generic map (
      C_BUS_WIDTH  => 2
    )
    port map(
      Clk_A_BUS_IN    =>  tx_TagMode,
      Clk_B           =>  AXI_STR_TXD_ACLK,
      Clk_B_Rst       =>  reset_tag,
      stable_for_sample => sample_axi_str_config,
      ClkBBusOut   =>  tagMode_cross
    );
  end generate;

  GEN_NO_TX_VLAN_TAG_CROSS : if C_TXVLAN_TAG = 0 generate
  begin
    tagMode_cross <= (others => '0');
  end generate;



--  TX_PAUSE_REG_DATA     <= tx_pause_reg_data_i;
--  pause_req <= tx_pause_request;
  --  Transmit Pause Frame Clock crossing
  --    Data must to stay in sync with request
  TX_PAUSE_FRAME_CROSS_I : bus_and_enable_clk_cross
  generic map (
    C_BUS_WIDTH  => 16
  )
  port map(
    ClkA          => bus2ip_clk_i,
    ClkA_EN       => '1',
    ClkARst       => reset2axi,
    ClkASignalIn  => tx_pause_request,
    ClkABusIn     => tx_pause_reg_data_i,
    ClkB          => tx_mac_aclk,
    ClkB_EN       => '1',
    ClkBRst       => reset2tx_client,
    ClkBSignalOut => pause_req,
    ClkBBusOut    => pause_val
  );

--  tx_ifg_delay         <= tx_ifg_delay_i;
  TX_IFGP_CROSS_I : bus_clk_cross
  generic map (
    C_BUS_WIDTH  => 8
  )
  port map(
    Clk_A_BUS_IN    =>  tx_ifg_delay_i,
    Clk_B           =>  tx_mac_aclk,
    Clk_B_Rst       =>  reset2tx_client,
    stable_for_sample => sample_tx_mac_config,
    ClkBBusOut   =>  tx_ifg_delay
  );


  TXCLCLK2AXICLK_ISR_1 : actv_hi_pulse_clk_cross
  port map    (
    ClkA               => tx_mac_aclk,
    ClkARst            => reset2tx_client,
    ClkASignalIn       => EMAC_CLIENT_AUTONEG_INT,
    ClkB               => bus2ip_clk_i,
    ClkBRst            => reset2axi,
    ClkBSignalOut      => EMAC_CLIENT_AUTONEG_INT_CROSS
  );


  TXCLCLK2AXICLK_ISR_5 : actv_hi_pulse_clk_cross
  port map    (
    ClkA               => tx_mac_aclk,
    ClkARst            => reset2tx_client,
    ClkASignalIn       => tx_cmplt,
    ClkB               => bus2ip_clk_i,
    ClkBRst            => reset2axi,
    ClkBSignalOut      => tx_cmplt_cross
  );


  RXCLCLK2AXICLK_ISR_6 : sync_block
  port map (
    clk        => bus2ip_clk_i,
    reset      => reset2axi,
    data_in    => EMAC_RX_DCM_LOCKED_INT,
    data_out   => EMAC_RX_DCM_LOCKED_CROSS
  );


  CLK2AXICLK_ISR_7 : sync_block
  port map (
    clk        => bus2ip_clk_i,
    reset      => reset2axi,
    data_in    => EMAC_RESET_DONE_INT,
    data_out   => EMAC_RESET_DONE_CROSS
  );


  TXCLCLK2AXICLK_ISR_8 : sync_block
  port map (
    clk        => bus2ip_clk_i,
    reset      => reset2axi,
    data_in    => phy_reset_cmplte_intr,
    data_out   => phy_reset_cmplte_intr_cross
  );



  GEN_TX_VLAN_TAG_BUS_CROSS : if C_TXVLAN_TAG = 1 generate
  begin
    TX_VLAN_TAG_CROSS_I : bus_clk_cross
    generic map (
      C_BUS_WIDTH  => 32
    )
    port map(
      Clk_A_BUS_IN    =>  ttag_reg_data,
      Clk_B           =>  AXI_STR_TXD_ACLK,
      Clk_B_Rst       =>  reset2axi_str_txd,
      stable_for_sample => sample_axi_str_config,
      ClkBBusOut   =>  newTagData_cross
    );
  end generate;

  GEN_NO_TX_VLAN_TAG_BUS_CROSS : if C_TXVLAN_TAG /= 1 generate
  begin
    newTagData_cross <= (others => '0');
  end generate;

  GEN_TX_VLAN_TPID_CROSS : if C_TXVLAN_STRP = 1 or C_TXVLAN_TAG = 1 or C_TXVLAN_TRAN = 1 generate
  begin
    TX_VLAN_TPID0_CROSS_I : bus_clk_cross
    generic map (
      C_BUS_WIDTH  => 16
    )
    port map(
      Clk_A_BUS_IN    =>  tpid0_reg_data(16 to 31),
      Clk_B           =>  AXI_STR_TXD_ACLK,
      Clk_B_Rst       =>  reset2axi_str_txd,
      stable_for_sample => sample_axi_str_config,
      ClkBBusOut   =>  tpid0_cross
    );

    TX_VLAN_TPID1_CROSS_I : bus_clk_cross
    generic map (
      C_BUS_WIDTH  => 16
    )
    port map(
      Clk_A_BUS_IN    =>  tpid0_reg_data(0 to 15),
      Clk_B           =>  AXI_STR_TXD_ACLK,
      Clk_B_Rst       =>  reset2axi_str_txd,
      stable_for_sample => sample_axi_str_config,
      ClkBBusOut   =>  tpid1_cross
    );

    TX_VLAN_TPID2_CROSS_I : bus_clk_cross
    generic map (
      C_BUS_WIDTH  => 16
    )
    port map(
      Clk_A_BUS_IN    =>  tpid1_reg_data(16 to 31),
      Clk_B           =>  AXI_STR_TXD_ACLK,
      Clk_B_Rst       =>  reset2axi_str_txd,
      stable_for_sample => sample_axi_str_config,
      ClkBBusOut   =>  tpid2_cross
    );

    TX_VLAN_TPID3_CROSS_I : bus_clk_cross
    generic map (
      C_BUS_WIDTH  => 16
    )
    port map(
      Clk_A_BUS_IN    =>  tpid1_reg_data(0 to 15),
      Clk_B           =>  AXI_STR_TXD_ACLK,
      Clk_B_Rst       =>  reset2axi_str_txd,
      stable_for_sample => sample_axi_str_config,
      ClkBBusOut   =>  tpid3_cross
    );
  end generate;

  GEN_NO_TX_VLAN_TPID_CROSS : if not (C_TXVLAN_STRP = 1 or C_TXVLAN_TAG = 1 or C_TXVLAN_TRAN = 1) generate
  begin
    tpid0_cross <= (others => '0');
    tpid1_cross <= (others => '0');
    tpid2_cross <= (others => '0');
    tpid3_cross <= (others => '0');
  end generate;

  AXITX_2_TXCLIENT_FSM_GO : actv_hi_reset_clk_cross
  port map    (
    ClkA               => AXI_STR_TXC_ACLK,     --: in  std_logic;
    ClkAEN             => '1',                  --: in  std_logic;
    ClkARst            => tx_init_in_prog,      --: in  std_logic;
    ClkAOutOfClkBRst   => open,                 --: out std_logic;
    ClkACombinedRstOut => open,                 --: out std_logic;
    ClkB               => tx_mac_aclk,        --: in  std_logic;
    ClkBEN             => '1', --TX_CLIENT_CLK_ENBL,   --: in  std_logic;
    ClkBRst            => reset2tx_client,      --: in  std_logic;
    ClkBOutOfClkARst   => open,                 --: out std_logic;
    ClkBCombinedRstOut => tx_init_in_prog_cross --: out std_logic
  );



----------------------------------------------------------------------------
--  Tx Interface Clock Crossing - End
----------------------------------------------------------------------------

  --------------------------------------------------------------------------
  -- Instantiate receive interface
  --------------------------------------------------------------------------
  RCV_INTFCE_I : rx_if
  generic map (
    C_FAMILY                  => C_FAMILY,
    C_HAS_SGMII               => C_HAS_SGMII,
    C_RXCSUM                  => C_RXCSUM,
    C_RXMEM                   => C_RXMEM,
    C_RXVLAN_TRAN             => C_RXVLAN_TRAN,
    C_RXVLAN_TAG              => C_RXVLAN_TAG,
    C_ENABLE_1588             => C_ENABLE_1588,    
    C_RXVLAN_STRP             => C_RXVLAN_STRP,
    C_MCAST_EXTEND            => C_MCAST_EXTEND
  )
  port map(
    RX_FRAME_RECEIVED_INTRPT        => rxclclk_frame_received_intrpt,
    RX_FRAME_REJECTED_INTRPT        => rxclclk_frame_rejected_intrpt,
    RX_BUFFER_MEM_OVERFLOW_INTRPT   => rxclclk_buffer_mem_overflow_intrpt,

    AXI_STR_RXD_ACLK                =>  AXI_STR_RXD_ACLK,
    AXI_STR_RXD_VALID               =>  AXI_STR_RXD_VALID,
    AXI_STR_RXD_READY               =>  AXI_STR_RXD_READY,
    AXI_STR_RXD_LAST                =>  AXI_STR_RXD_LAST,
    AXI_STR_RXD_STRB                =>  AXI_STR_RXD_KEEP,
    AXI_STR_RXD_DATA                =>  AXI_STR_RXD_DATA,
    RESET2AXI_STR_RXD               =>  reset2axi_str_rxd,

    AXI_STR_RXS_ACLK                =>  AXI_STR_RXS_ACLK,
    AXI_STR_RXS_VALID               =>  AXI_STR_RXS_VALID,
    AXI_STR_RXS_READY               =>  AXI_STR_RXS_READY,
    AXI_STR_RXS_LAST                =>  AXI_STR_RXS_LAST,
    AXI_STR_RXS_STRB                =>  AXI_STR_RXS_KEEP,
    AXI_STR_RXS_DATA                =>  AXI_STR_RXS_DATA,
    RESET2AXI_STR_RXS               =>  reset2axi_str_rxs,


    RX_CLK_ENABLE_IN                =>  RX_CLK_ENABLE_IN,
    rx_statistics_vector            =>  rx_statistics_vector,
    rx_statistics_valid             =>  rx_statistics_valid,
    rxspeedis10100                  =>  speed_is_10_100,

    rx_mac_aclk                     =>  rx_mac_aclk,
    rx_reset                        =>  rx_reset,
    rx_axis_mac_tdata               =>  rx_axis_mac_tdata,
    rx_axis_mac_tvalid              =>  rx_axis_mac_tvalid,
    rx_axis_mac_tlast               =>  rx_axis_mac_tlast,
    rx_axis_mac_tuser               =>  rx_axis_mac_tuser,

    RX_CL_CLK_RX_TAG_REG_DATA       =>  rx_cl_clk_rx_tag_reg_data,
    RX_CL_CLK_TPID0_REG_DATA        =>  rx_cl_clk_tpid0_reg_data,
    RX_CL_CLK_TPID1_REG_DATA        =>  rx_cl_clk_tpid1_reg_data,
    RX_CL_CLK_UAWL_REG_DATA         =>  rx_cl_clk_uawl_reg_data,
    RX_CL_CLK_UAWU_REG_DATA         =>  rx_cl_clk_uawu_reg_data,

    RX_CL_CLK_MCAST_ADDR            =>  rx_cl_clk_mcast_addr,
    RX_CL_CLK_MCAST_EN              =>  rx_cl_clk_mcast_en,
    RX_CL_CLK_MCAST_RD_DATA         =>  rx_cl_clk_mcast_rd_data,

    RX_CL_CLK_VLAN_ADDR             =>  rx_cl_clk_vlan_addr,
    RX_CL_CLK_VLAN_RD_DATA          =>  rx_cl_clk_vlan_rd_data,
    RX_CL_CLK_VLAN_BRAM_EN_A        =>  rx_cl_clk_vlan_bram_en_a,

    RX_CL_CLK_BAD_FRAME_ENBL        =>  rx_cl_clk_bad_frame_enbl,
    RX_CL_CLK_EMULTI_FLTR_ENBL      =>  rx_cl_clk_emulti_fltr_enbl,
    RX_CL_CLK_NEW_FNC_ENBL          =>  rx_cl_clk_new_fnc_enbl,
    RX_CL_CLK_BRDCAST_REJ           =>  rx_cl_clk_brdcast_rej,
    RX_CL_CLK_MULCAST_REJ           =>  rx_cl_clk_mulcast_rej,
    RX_CL_CLK_VSTRP_MODE            =>  rx_cl_clk_vstrp_mode,
    RX_CL_CLK_VTAG_MODE             =>  rx_cl_clk_vtag_mode
  );


  --------------------------------------------------------------------------
  -- Instantiate receive interface
  --------------------------------------------------------------------------
  TX_INTFCE_I : tx_if
  generic map (
    C_FAMILY                  => C_FAMILY,
    C_HALFDUP                 => C_HALFDUP,
    C_SPEED_2P5               => C_SPEED_2P5,
    C_TXCSUM                  => C_TXCSUM,
    C_TXMEM                   => C_TXMEM,
    C_ENABLE_1588             => C_ENABLE_1588,
    C_TXVLAN_TRAN             => C_TXVLAN_TRAN,
    C_TXVLAN_TAG              => C_TXVLAN_TAG,
    C_TXVLAN_STRP             => C_TXVLAN_STRP,
    C_S_AXI_ADDR_WIDTH        => C_S_AXI_ADDR_WIDTH,
    C_S_AXI_DATA_WIDTH        => C_S_AXI_DATA_WIDTH
  )
  port map(
    -- AXI Stream Data signals
    AXI_STR_TXD_ACLK                 => AXI_STR_TXD_ACLK,
    reset2axi_str_txd                => reset2axi_str_txd, -- from reset_combiner
    AXI_STR_TXD_TVALID               => AXI_STR_TXD_TVALID,
    AXI_STR_TXD_TREADY               => AXI_STR_TXD_TREADY,
    AXI_STR_TXD_TLAST                => AXI_STR_TXD_TLAST,
    AXI_STR_TXD_TSTRB                => AXI_STR_TXD_TKEEP,
    AXI_STR_TXD_TDATA                => AXI_STR_TXD_TDATA,
    -- AXI Stream Control signals
    AXI_STR_TXC_ACLK                 => AXI_STR_TXC_ACLK,
    reset2axi_str_txc                => reset2axi_str_txc, -- from reset_combiner
    AXI_STR_TXC_TVALID               => AXI_STR_TXC_TVALID,
    AXI_STR_TXC_TREADY               => AXI_STR_TXC_TREADY,
    AXI_STR_TXC_TLAST                => AXI_STR_TXC_TLAST,
    AXI_STR_TXC_TSTRB                => AXI_STR_TXC_TKEEP,
    AXI_STR_TXC_TDATA                => AXI_STR_TXC_TDATA,

    tx_vlan_bram_addr                => axiStrTxDClk_vlan_addr,         -- : out std_logic_vector(11 downto 0);
    tx_vlan_bram_din                 => axiStrTxDClk_vlan_rd_data,      -- : in  std_logic_vector(13 downto 0);
    tx_vlan_bram_en                  => axiStrTxDClk_vlan_bram_en_a,    -- : out std_logic;

    enable_newFncEn                  => enable_newFncEn,             -- : out std_logic; --Only perform VLAN when the FLAG = 0xA
    transMode_cross                  => transMode_cross,              -- : in  std_logic;
    tagMode_cross                    => tagMode_cross,               -- : in  std_logic_vector( 1 downto 0);
    strpMode_cross                   => strpMode_cross,              -- : in  std_logic_vector( 1 downto 0);
                                                                     --
    tpid0_cross                      => tpid0_cross,                 -- : in  std_logic_vector(15 downto 0);
    tpid1_cross                      => tpid1_cross,                 -- : in  std_logic_vector(15 downto 0);
    tpid2_cross                      => tpid2_cross,                 -- : in  std_logic_vector(15 downto 0);
    tpid3_cross                      => tpid3_cross,                 -- : in  std_logic_vector(15 downto 0);
                                                                     --
    newTagData_cross                 => newTagData_cross,            -- : in  std_logic_vector(31 downto 0)

    tx_init_in_prog                  => tx_init_in_prog,
    tx_init_in_prog_cross            => tx_init_in_prog_cross,

    -- Transmit Client Interface Signals

    tx_mac_aclk                      => tx_mac_aclk,          --: in  std_logic;
    tx_reset                         => tx_reset,             --: in  std_logic;
    tx_axis_mac_tdata                => tx_axis_mac_tdata,    --: out std_logic_vector(7 downto 0);
    tx_axis_mac_tvalid               => tx_axis_mac_tvalid,   --: out std_logic;
    tx_axis_mac_tlast                => tx_axis_mac_tlast,    --: out std_logic;
    tx_axis_mac_tuser                => tx_axis_mac_tuser(0),    --: out std_logic;
    tx_axis_mac_tready               => tx_axis_mac_tready,   --: in  std_logic;
    tx_collision                     => '0' , -- half duplex not supported. tx_collision,         --: in  std_logic;
    tx_retransmit                    => '0' , -- half duplex not supported. tx_retransmit,        --: in  std_logic;

    tx_client_10_100                 => speed_is_10_100,     --: in  std_logic;
    tx_cmplt                         => tx_cmplt
  );


    mdio_i_temac <=  mdio_i_top  and (mdio_o_pcspma or mdio_t_pcspma);

    mdio_o_passthrough <=  mdio_o_temac;
    mdio_t_passthrough <=  mdio_t_temac;
    mdc_passthrough <=  mdc_temac;

    mdio_o_top <=  mdio_o_passthrough;
    mdio_t_top <=  mdio_t_passthrough;
    mdc_top <=  mdc_passthrough;

end imp;


